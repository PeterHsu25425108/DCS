//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
B+IIvQa8RX9wPAaypmU/V4zKifoT46r6vphWfKTKTP8WS9AQmzlm7OF6ZT9kO3o2
ybocot+N+YyO0DGJw/NAnK4or+tZe7TBdZZXfgZG4lHnT0xzH1BYa6HympkcJmfP
g6gEKm8omk2pUxU2R7fbo8U6Pn9+pHIZV5s8vSTtX7BJm1Q/K1b796VYGync2bgl
hT9x/UMbJr5fMcIas7j4pTQsmOLZ6JswltuCOS4ifSOplcyGzEg5fMbC7LVAU1jb
rFdCk2mmj05GXpI9WX+4T0bL1A6NvFHZLHw8GnFPhHX2Mpesqdf01FTmi02itDG2
IsG3L8s68IXBgKG9+RHYDQ==
//pragma protect end_key_block
//pragma protect digest_block
16ua/d8FEZS/B/Kh8+o0ejZZ2aM=
//pragma protect end_digest_block
//pragma protect data_block
p/iSL+u2RSHD2SddsMqZDvk/xb4wIaXpMC3X/c7KAjYDyyYP8gRuWYkcUn2Y19o2
K+fD2TFVsDoWLhspu0drv7ivlx+YfHb+AG5q/AX0nVvNqwSA13H7gKbdwGYe9t4J
GC1TH2ety/RIVfliFb+gj0MdyxEz3DU9WIaQi5HiebR3NWpneSjJyEvjnv/9CU5E
sNtU5aEgPd+ILdCOUJ1O3BQGANZr3QbK/+Ecv8HurNFedPpemi0AeVlQwOb3NCMG
Fok/nM/btI1vzwmu78RoBEUp17rQFoHKd7iowzMw0G8kBMLgu/EiTGkr3rk0Rd24
VaSkjXs2LVjJEcIhaJlWWG0elTicNB7HuKT81MeMozwXiE3uR/8FCin9WPQ4KFD2
VQiyQJifU//x3Rs3z0+twlPRo6wGUIT1A9q3lzfl2q8a4TLFbPTWAg+feXLYyvRA
3lVKjyrmpn7hOGOre90SXfrshBq6gedmrZJX6ZQkc8NAE2b9IH8bJGb89NXr58Jl
ciCJzK9WZ7BwHtF/7U0Zfh/oPmdrqCb2U6iTYXRNLCLWtSVGepnOM2Tqe/06/E7B
yghhnQ2lyGqYupD5w+Z0dKjVKVtCUfDSS589o040ClkV/Q9v1j33pcHzoEFA5Xs3
ny9pO/aATnpzLupUM19Ap7KGP+o/a375npKsOMfa6EfW5qRFkVU9cKeSv0Kj/D5/
3nOiDaSqjILdSUkvcq5XxbMM4YzK9n73hAz7jUEMXocTPOxK5M3nIsoLf9IVGZIy
9qnzuKePvhFmNQgQeSGKZn+bgztmMJ6WDyYmrwz96PveVOFEH5GaH5N/rn647DTL
LWVDaZb9u2b1v7eXJpCaCaOjr1JtWSKLvazYbbll5TXnaIkLS4ZNqlGmx5rEYV3j
c96dC4WiTHBP5fL7/UgpUIsAgh0i+93+s+JSZDIhm8QIZyI+cCMLqb82fb/V6Trw
DUUnpuWmprPPS/WMXWaBaUJDivA8C/nzoPNni3j0cM63HHc96nD6lLcpF4WRhFdq
0iXV1caXbbRwskFrQwimczKptFpkOFcMeSCcDsA8fg1E5mrfQqU9/y3DclriktTY
HtggJ2xVT0ru2B5M7XqxacoJi7ciY967owcjmmkDesAP20MYzBadsIcj//hCJMv1
Wmc8Pha3U8Dw4+56t4JErTUlIrdjcfb3YUtegRg2eG3tErkkn6rMzF3q1+avAOyJ
ipGar8l0ZgNx+xEN11Kn5iPzj1mcfWPHZMRoEF0nT4iUtvK+ilS2JMnhLbNps9Vg
u320kKGeX/bG9tUMeEPC3eUkaGMSWb2zhMJ7hLEPX52bppseYjzx4aSdleVIBBGm
ETQs60Mzanxaqv1sbAq8Gytm2njtnYdwdAhAODWjCP2eAe6RH4koPzWnpizbuvmU
Qo9KFwxKTjtWlatfi+jby6HvdoruPQa6XKIRN1VUOCYD0ijuqlb5qBuuKMT1ZkEp
WIEj8RtwisMqFHXrNi6Ry9969x5elHHFjufQQxlZKLqZQZKyViDPgPwQpqd7F4FQ
lFXB5SINjtCkxFOU0LPFyWtkZsuFVtlEWbPJrpnuApx4T7bVxeLfpWYQhfe+1HoD
EMBkUWVH5oOL/OxdQe94Sy03RJ3TT+LGo3/ecaVmt2+UwCaVfA7i2Yfzl+38TNoX
2urowqOHiAkgihz0teEYK+e+giSDYvIzt5TYO2dser9xdSmHwTDILGcZ7/Qsva7Z
ZXfEgjY4l/LsqTVx5jzLD/X/Jcc3D2uw9FDKGBUXjJM1nMEmrpoVWDnzrdTdFTJP
sGfk1rGsL+6We9QHA37htv0x2K9CEJB/NxaVNENKR+tjI+hePYS+a+CsNo51S3g2
Ia6Na7uag2slKwQ7BPXZyzDh1OI/aR6vn+pTMy9cWQTpaLdtCDd3INW52jzt7FGT
gwWnU7XnbxYJwTNENvIVdjoFfRrxdXNdENptdhxwoW2PR5CCz1WzMXBmraqCPwfn
39b2buZVZm2hcKSYULVBMyHspTJ6k/5aHY8I4OKE5q5jd6Z1zejOSfgUjSzKKaiJ
e9zAhMxxnldYRdfh09BwumXbYKYwIONilScAOqZolsi9ejNzJjw+C/IxE/xH8kT1
m3oV8wH7Fv/cla6daIZ6Pnre64ouFbpwwGXAl3lB0W7OoNl2wKInlQVLSWWTCVT0
YDc6PEqqkIn4Idvh2aP2yzmgEGR4Hb3hq5MdGAJgYNZdZbxsM4dlAoWXcTZxazrT
69EW4kb8j7IK//XMNtMc00qNWDLj2wWxJRmVrYPHunBYzpTOzcmvNM5orsJQx1kM
JaGGNGMpVCUuL9mta6WEZv1tsQlhIzlUK6oRMkvcoYVS5nxQ8mEXT84WWhqtXy8I
JSRTJldyyqiB4f4wZWGRxPA4eqFMsJltHb3FYzfO7APxgMj4iq9Ikmv4djdnGuMS
gPm12UxLpf84UFBMoTEGakXN9AMNgEcGj8ygfG10okgWa7NDvkNoV5k4hsOegXWE
3oi2/iizvElXRgG1zUq2BcaU5SA5sWjWcPbTwn+2RVMTKQdKwu8nzZOhS/cVtLa/
pEXy5J4Y13I1rkr4dr85bo4xrFY1NIWfJeSVH+esNWsBVgaldwjlkP7NhczKTycl
u0Fp2+WdmH5FKwmV3Yi0NXl+K0d8ShqUEmPvlWsh/PnRbnwzPLVBMs+0YugOKUTq
9GeQ/wORVnaTplNfXj6uaV9Hu/UHkfEleW2jMUQw2d1MYwt5qGO6pDqhuhsRifmS
zt1OOQuF2FFH4a5g1tUzMa8Yst62jftxb760R2He68UFWD/hWxCN5F7fiKxwlnaZ
Jexo5jY6Xm3s0GF9C3sWlebGNumSmtMdZr/FVvzkDva8pKOdaS3y2MlNbAFhV9Ea
kKb85zWNyB12xRThPSHYFwcioxFdph5MKKTSRvcL18SyUv8ckbz0pFpEnurJKSZs
6SlAAaT8NIChonG5B/byKFY589U79awUXZKI+K1t0Vv9SxRXSWhz/ImWSNVh8s4r
xAMAO0QD/07xviaOaXN7EgPRSzHbU8On/XOcEGdsVwATus3k1QgHDp6OcTvccyAT
rBMWmJYomUlIrawuAkHrAnhXHh8xj5Q4PtCsKbxmv15WNd3TgD0inFkTQ8As2XLk
+G+x9ezrgM37mnMKqv1QaP0noXO1h6QYEsrTwLlXLAWUiX9LHmpv/RmNPxWv/IJz
17dEVA5TGepNEU807GyXd/6ZnXDSo+04qHLjHxurUkoQQaFWuPeR5EaXYGbMDsBo
g1iG43qHa2Uvvx3vygnbvZDuQd8dwDLBqWTPxn4cLu/wFVpWf+N3Ku/1KJEjyZbX
sxk0Cx4bmMN0YNOGVyKZOfhfliDdlgSvwtMu280j93c9cCUKIBZr0k9jGDg9p+Ot
WvrY07YtWEXlH37AO5Vo5ZD3Yt/+BozVbwz0+0/h8Q6FtE6iS+ei5dPL7u7PgdB1
nk8OeCZxfEd7aukAUn1TawhKJNOu3P8r0wKn53TkclW7MvqWw7JgtgCITBUiUXcy
dEd7n2C949x2u8oZROPXTJEsG1wqD5xHp239konAAeknFdLOJYdZNZZ3mTEK0vaY
shCIfgbDTj8clUu2p0XZWZbZz1reYSexdDuyq7Og8e1I3mnNo+kww6I77nEOoD9R
0KaidT4VLHojMqlLBBZ7d6+6/5tarV1iwPSjXaQi55LNFz5ESfVFJb1TUiVrKt+o
BYOKDtiO96ySqWQW+R9FZbr0CGOKvPyGrMwUWe/1fAn4OSrSabw/sDCMzAsuF0wZ
mGfMuibzrasFmCyl+LfwZhczEQoIryovczXikT1NqxhfUV9aFmYsseRgEJOXEw6D
sr4VjmyYtX/LTjBpVu255LCIXpGX39zApB5FRAmYgfp/9lMN/4IjZPyFavBsc8d4
DovtSh4L+93QV+4loIA/V7v8u8nFQD6/2pfe0JhvgcLpyeApYrqsEkoadGnSkODo
UDuYYSsieBa09oyOvKnIKNV0Y94Y3UZhJqGcCD3Y6dir0ZiyN+AC62JjJwQZtVV6
GnfudWwr8xpEhsAqBAqUra/zhXGJsYhscLnjsl9Y/DmiO+LxlRdt+3WFiQAdidt3
WeqjnsEtmsOQDPLEYAVq+91exNIHm6N7tV5bZA00gCj+87iQGN38cWe/z2Ebvh5J
WZpgyeMQCHP7quLoCVUfyqDbux119rl5VMGo7rNqQi032YB4Tur4qmoUwyCxJpo6
Owj9nLVqui5rtvtM49tKnWQBbEQDW+V5YoW5u5zGwgGh9eZvtP8wfcW8yCsLeB68
cfndfjxn0wF6OR+kOp84e6d3iPYy8geF9lvFksseEQ7Lvdx/faJBb3vu+WvExKkW
/A0tNWUwfLei8GG6dB3MfWugMGfC2y0FZU002vEesYMUkWBHqiVXZ+5GnipaeE73
fsvaMm2JnADQfyA8DYQlx07S9IhPMIWh0GGOGzkSG4AXo1oQbn+Q7nkTKJZYCPot
e/w2g8i5AzYVfjgExcqEnJGP9H4Kzshib+jtOEYjmlp6YFtPWtmTtKvzsBw/SCuq
KmXH9jcj4bAnGDS+yFlXBBtD4G9qVVbWAB9WDnxNJFaqHdyLOypvdPCcVTYHNhjH
57FN512/1MD0Ls4kaxOlcQpj5YVdViBarqqZRvgynRpt/vNHTQziY8FVzKK6VYyn
FQuGtScW+V5Txqhu14EXRtwhEB4FjB9YN2+15QrLUj6ohG39swJTZOkxmDCvyphE
iS3wWZNF2gtYZeAfouO4QhlX9UqcFV5ubWvC7Aibyz6nUXMi0eUbp9RecCEn4PVE
1o/gUXRxfAosymcicDd3a7T8Bh9dzRaHnokobcM2OdNiBAPZRu93W7ePrExr/zFx
UMKvr/9grEq9W14gIt+BTbFntS9yULHE/Nkr2gVNZu8BPT46VQSAEvMDPXtHyDWz
bviX7xzJ++6OZ59GxLgZUfY6qiaQhPs9tzNr5Xk+qDq464GuFQ/lZt1nNw75KI1U
vF6/5nFr4euvJ81KBh4+NOfygk9hg7JIowLvWbhsjnE2/mCi1Vlv+40ya590+Nmy
aU9Rx2VPieSvU0TPydzTcj0Kuw10bKnnu72Wc3YvrQQVaZ8V9T9Pkk3DzoQ1nMiB
mZEvzFhGAfg+GZt8y7IzpzxsbkIhfJOiQs7cubSM16tpzUiW+1gSkKo2Da+0AqW4
9Mrm+JFfM77jGUJEXI025Vn5RIOrR5YebltdwWbE88pih4vMBbwEHeuJbLjaAIG5
ko6lJ9qYhVl+QRSmTPdfZR2YPGc5VcbwT2fKLZF7wID2HVXo7semVl87JJgJLevs
ZYsL6VmqScfD5NimQ3iRvtNpom/l3Djh6qFDWb7B7+b0OGu9btEzqzgIqENTE+tU
ib6Hke6SW5Ee02NUTOcGdIkzZibKyEQbrPAsp8GKWT67Qwvo3xMjYWz2/Uy8Uav7
xFmk71f8XJPZu2yG8+MBe6Q+q/eHPjfwNfTgCrDTRfXAXqgwe/jxwEkiJiDXDtg3
rWZDPx2sJxgPnuGLAlODbhLxnbxx8J5T6uuaku+CcwsTut4ekEH3xvQVMOIiayHw
w+tg9JlVkjanx3NdMVHGFATj70OKsQ01XSt9PaEyx31qs7jSjiziKoeF63ub0M+K
j16BiLW3uPGj3czKkate+zafCitajjUlG6rLW5QOzQcvNb662x5T8dg9CcD+sc5H
W88wxbG/NrNpnjcSZsWxnu/74LU9yV14M49RgwHmR0yzdpP2kTdz+ZSR+3PMm5Gl
wsM5svzN2XUeTTQ86BtAUHVs4armEOSCfvVHMEWkeA3oXuV0HNUclKLdKpkIm0Sr
hQGvBMWPWT1bfFYN9oEUPNPFTFPKNhz2os+JYyVcnXwHE/tbVqP6FYAkau2RogqA
ZqMN/AejLQonbmLaiHEqWfHFrqFsr8IlX73Lo0mJhbmtZ1RMEHVARNi+3yp3AXJ6
6VuFzzIs/CoYtKBVwP9xnIxrJgywUNYnx7e7W1atVKyq+yMHSMvk1ibs3IKwNQT5
8lvzC5xkBDE3ff6SLqS2vXaHJ971Z9AJkYDwqR1G1K+kD5g/GkWqvvjz1/QYK4lm
V4KViqoCFQzyxyf7Y/ktTCrx7VozeHQ2J1UhCrBD07CjTPLRSLvjgB/VR9YrtdzB
WVn1SEYjCPxLHBizy9/DeqCF/WBGwO/lx30VDdsL+26ieIOFyXVZYxrW1/beWBah
bDTQLespkVvvDueUK+/yBKYZOahta8RE8hxi4PdE2iyd+VZvMasFDFwttnk3/Vx4
G7VzC8rCWEfZB6NLYKhk2IK787HCPzDd7tu8hTlN3zON3LM50gWzS6Wn1/RZJlWV
XkJHZDzvmkdGC9xxmoc7rCot67dLuOLkseubA0J95sZFY+IUViBTba3Mt9Hz+Evg
G48o4UQPbkWhY7LhtoX6BLR+OCeg+964T7h6bZdMWNRUkQyrbjPsjYnZbG4iwxOe
6G7dxGzDl97JoGTWc3gZdsfuAcMp7W4QFXGQ7g7UavSkJ6T2IXQ8qFkSj5+EpULq
sL1h8DMJ7ZJHtmBXqGQh2h4NX0cO/dKMyJMPdVAoVShLKRaiM8f88s3DuiulLoHp
btxXSGEkyb/Dhylvs0xDobBVwmurg0PNoK4eXlVBMyqGkOQlCxA+k/sNzkl99SEK
LKB7xX6D56hjav9CIsaDaDPGTnJsxz/u6RpnyJ0Y1SbTUCPKdrBOx4vh5/KjZ1kK
e9YKLr/Wg30hmIidYT38AX41s5ZQIbLO7Nu3MhaJ9YruffUd1QNZzG3jZesZk1+U
k98FWRDKZ+UGU6cIp11JZyeMwNR9Tt2wJRdpll63DjxUwcYKfpRkJfizY+oUIBsD
warGJoe59RaP+7zktZR36aeGXJMTzoxz8i16qkDt3IzDnrbKMFnTS7tn7rcpQM1A
Glsw8RaOBM+3FcE3UkLYrmmaGOpX1eoQVR/6eXFxFlDsYJXNuIlSVKkdk1VaNWEC
V8TX48WH0e0mQ1HB4CSI+0jdGkoaK7qhcKDFBnLibKrfF68cNLbtOdbzPblvcDvU
AqoBGSLrzrtcbz/Qbl00IlGLsVutylPZXJqslauqPYFBvO4/GriKcfweNQFuNIbG
uF/jh/Qnb35f00Gs+OczEM06uvaxzVNfpQq4lLZxp1PjjxIsz+PLNXzijxulgzzU
ux1/yiAQuVnbEDBUgW/JKb4vofaV1eSuMvWBPa2B95JTXTZCLfnpVXrorYGajUwJ
pcIwHx4yL8CsWBcrCKhLrmTK2+j3eo16A4FkL5+MWgfiUFnBtHmyahRuVpqt3YcR
mCiKXpELIjkvfUw0tUKVKPfNZsukWt4E+T/L1AhU14NnmADw/8JgogT5L8SEQOQx
yBOt7tOa1OelQFrk7fcloaPlMTtZB9SEKuxXJ8YYghCgebdDzrNN4VLb/ukuWHM1
Ffqlj8iII2nYAvADHtIuB343lhNyY5cakXo/y4qMai2Kgn5f9A4aCPF5GZadbHk8
R9hLsz1CN/O+w+fzijl4gKk+bePh8tsiUg4oI6ofMIYiYZMHBaL9Ut//+Q0Ei1MX
C+1GSGNqiArhZ0KS5kF8LhI7UEuUyQ2rrCOwSsQ45q+EKsFPGeFp01Z81FuagnXQ
0EUrJ6UudWdeaObnwKhIixefnqNe/Ub/eVuNGI9SbMTyT4fhKgCmUi6D6ONpn6/n
Z8hWf1zF4/RI8lvNdh0Fsvp8nIMup+XFClUclCt3znU6qR63ZKbg6qWepZj81rB0
WmE1qX1AVWESjZjVvUpIlnaK5BUpGwYOkToNBGiFl7edSBTuo8Qljzgf2pyWW9xj
DIZLL00HKvBxurHFXQWRQ2tbDIJSJo42/Ge6ahkf1m7jtR6aoj9YG6WrdHjbxruG
4BWWt9leMbKSN245TFK9AeET+Elfn06r8zb+cWVTtrHaYEOovnXdTSsPT6jwNLnt
SkGQbITc18sq7AFrBYhlJ0li+WMGCmJz4FJxdt5nL0aDo7qcMJi/3cyflkpFd8rs
7hv2JjXRGdF8NIRVrA5PCgc+P+u4XuMANPg5UhxQa/DsUH1e3CjEXN3TXK3qOTUD
8fX4Fi4QwqB57xFcqRfy+OhDCWNq+iiK5jVEczknz5t/M6hsT9qCE/N8TkzZhdBf
jJn2z4ju8oZhtKwUDYlCiPRipAPugeARJA/e1y1Jsrh+aTAByfoc4H2v6uKaz7DM
pHdkSl6D9EfvOcuY2gML9lxDBKePWwRDNZVWZUQuIncIXpiKmFMumc/cpEJhbMNF
yCPBnm5tj83FYabZQaTwAL6eJIMJIY3ZurZNoPEQKqZBoqcQERGwy4X0RAy5RBSP
ZQtjUSqR2aLRIBxU63PKYz4v/D/skPye0KqVw28sp8gcszURd9jWaPwOnbu/KkiZ
KNHiRlUYezcG1iGuhCL8ynBbR23Jiafz5onSqehI/m4YXZDN5uVEaA3DBkL1Bjw/
eyIOKacaSJZwsE1ZiFGjPXuwkkvBnC7gZmIpl9OitLCmB7pVz5jfSIo1dCYmTbEH
TID8yD7QlDa3z8i/zE9ZrvxAWMTB7TGjNFCE59w2xZAenXghhN+0shXFJn/8m4vZ
7C0mdS1f1w6bZQYy47frjh/BIAhjeu07uJi/amg0fxd1sXo+LRhx+hzst5buoaKu
QAHNW6ljKoxE77KLz6EPbA2Mql+VxDiTqwzo08Fkn5o95W/DTDi5QF48DPo/EC59
BwufzNLSGM3Xd9/RvK3mvkxZwzAYz+3ztCd3IZPEkiIGXAnlT181E5BQfW0GfCqQ
u/tL1DnC20p6aCS9HqRUa7sfQAb5ClPbfwEjXRyQ8cIytvLXNOLPAI8AOVvfnt3d
M2x/3r2DvcqZFzT4b4CWY2scbZ/AOs24XU1lKD9i5rvrBaJ+SjxB+n1+wgzuWUo4
0/vPjjoq1E6xEOdr2PyxMRUwKKFI/HqtC3vS6LSKTYFE31nd4+ny1cD/HzxdFFj0
tn+RSt20E2pPkvOi51Z8cNp0BBhtsyR4v0glDQ3SO5scZ+n+1RbbVWVXp34Q02M1
tlfR8xovAY8IslKdEZfj0FdH3ipdNC4WnLIzzOknT5PXeTLp/5zDjw8AOKhL7oeh
drHxEjvqgz0Eqj7YoTZ26dx5ZEBBnab12vI6czuVxHxhzMP8VQBO5yxyW5+0IvAm
7QmHF9t89Itnu+36ZyNYMCGoRHncAExcM4BzenoPPQsraCcM0bhvnF6lH7fkMjKI
lAi2U/a9gEIihIWT2knWWZUoiIvOR4t0zIzMfXMYx+H3HfxclKmcg0upVDvH42oL
yevFwDklUbmK4kGZdQwGt1hXAblSwpshUjN25qYKaFHBThKLAg/4g+3Cv+4Ug1Hj
uRb4ZGtIXTMxMkNUzl/JqG2lcZbycL8rxCP/rTxMUusrHRVvt5TGvPCqSto1sb/u
reRpmidwzGo22FghovzabOP7SLjdwP9SuvtKUwNdBRSg2VL1BZKQbUOjSEDkZ2fB
0IdMBHMRgo/WoQYo50kTvcVEH9jmx2wckEmKT8Sbr7AGyPazDdWTaziulBIuY+w3
5Byc5XXEw5pm0vt6FVl0QvIXx1uST0Wh9oKt7czGd7KtnG/pP+/f/K/eg1Q4zqLP
uMQ/fsAgPIkoTbv8qXxy/EUemF5K9mUjsZZM94AYq91zoQ+wcbnSD9RBq04qj2uE
ZTfMWCaXbRj//vblyXTNsA7a5Nx4fHt0llNIJkIOKIxxuiaShZX9J6kguArKE2qf
9FP/yyxl24oV8FmwWhqWulDMUTJ2K04hGa8ucbLXqnYgRbCNG5y26fGipkju++O+
tJSd+l61aNGaKPUnGggUAnwihjYi6SM6CuqCZ23iwEk5sXv6SOH88OcWj26w64YC
1WxEor1U8zxCO99UeT9Hhu9MtWlvB9yDLieej8UjTu6+H978zi50wzH2qMQYeA9d
WBTfcI5AYyJHUdS2GqjcyH74WzJuEJ6hnmsJEEp5RLb/9F/MQsBS+yyfC6b9IwwV
f4XLvwcOk8uZTjwa+44p720JrqrfOQIqK9c1K5tNDpgzvnOLUAqlf28niO3dUEnT
jZ/xn2zFGSfycURO64FgZ4HExoLV7xC4jf41i/q2QpnSXYmWSWishT3nq2zvWGy4
Ef1TQNtTubpgCNx/j6vqT3vA6l27gmzWVY6iRhZ1t5syowcFiZAnUGvUsWatGR28
yG/6LSopko34gHkdGZlShC2DRZ1wBXt8Pyp55dFC7a3G24GPNFftt7O6C52/EhtV
ZDRhJDhV1RALeDIo23l48zWe2rX5T7HLkFO9rVbHE443BN0Qum9DETffCszRdn8O
GaY93m01VTj0hGLo9ipAPFXaFe9FPuRajimrdyzY5urRWn/hQ319f8/zCW2o7jnJ
fTxkC2+Yq9bIG7Xajc/F0efYDL4rTYoKA8sfQhOpriigAR2yt1tXIxSC+R4P7+gr
mS96Mjzm4IVo04nQkt0fr27vkO8Yp2oGvrrXQrZ2eRwl4UIAsBwS+h2GA/EOHtk0
7TBi2B30rLv6qQwIGO5CG6l5O8bkPVoenHatmjBc9f2+XTBWn6urqsQQc7cj+qdn
9ml7Dz26tKMOzK4pgop5zQXttp6r8+4y6XQUZzOUzSfQ73Gb7QrI/klA5+5ZbuXD
iL04o4OdMtu4IeQnx19c9fJWzCmOetTXjfwYZf8a0KxrZoDHOCYyLbbCUgiisKIr
ndVMPdTEDtjlXOLAB5uq8SrGH+OlfGsylc41zZZLfPFSy4na2E2Wrdbxc2P9HrJP
STsdOMKvbRd1hR8oIXhsv6Z9AY4KKD2IWeteNyAildBcKTXFV961Rg5l3reqACKj
uE+pkkrmUUhonmfFdGCP4wvh4JqJtaWkB3yvwkGpIn8cGAT1m4tdPGLWiQsYUjBZ
vmgf0OlZlWLwRNy4P0qDgJvsF9k3IccwgbbLQRjL4gx9AszMu/FDQjSz4GIBZlhB
rkaM+084FuhxHHQrfPaYudlKqM/y5cfjKIFTi2NmFtaXmoeixAIDL5yuBoSfMEyO
YrE4/dlerjfRnaqM7aJL23dOrFo0FEBfjn5tBOg8cbAyVauxewHf6ZanWfCXCdYe
CF+lwcKvybwTFn3p3GxdniO5ntVlus3PFN9aWVehpdqPc7U5KVAIiikfD1DUvcf0
MPPbTgRvNBfc/zdtFxw1vtvv4UIlkGHp/KgyugoKnxP+6jBppe8A/2Smw/KJ6usA
ORqGc6ary2WwJmyyU4ICsck669/dzLDRvIiH0SZsbIz5G4CffgxaYVgO4r3Vvfln
CEkrgtmbnTgBvaH4/o4P+pv+lhy/6VdeDMstvUbfx1oBTOp7HLzydYIfMoUHcFdQ
c7gN4hwN+8hUSIEuHq5TbSYI18lr5zROvP4CUR6jS5tivIeFBG6ZRNcOejY3/641
cNoR8aB0jH+HRsnEQNZt8A6B9hXB+6lEp3unBa26X2dVoNx7Bm2A1A19y+CH4/Pg
DW6SOh9YeZA+Ab1Pj0PShZ6Eb7VMmq50b6z0LDx+6wNlbjQC7qYLoy0Evq/z0gpr
CTFHgmXpaxvpcuHIdDjr3oS1Lrp58GIQJqSfYXiX/xmvZSSA8w7odJhWdOMqe3uB
gOE9S2VV9ObrP+tmtA0UGftAEZ1xa7/dwMxjPEMYRJaLUGYj9pJEQB8Ih7pcOeAq
r1X60gGvUeKNip31wEqfgKxG9f4I+qPeWuOerU7nKxqGxrxweN2FWr+RWK8lhBrR
McRLcVvO0R+uD4skxkwDtGkKfdW4WgsQ2FfteBYB4uF4EC7EYGRzj4EVvuKF7LqG
4gmOoyUDSPkvJ8zvGuE+7kmg3nH8Wpy9Z90w1laFjM82YwT4bp6TwjTsl42rRw0R
9RmjW5nllW0WyzLO5lcMHss1VZa72TLJPT7sl7F+FJ8bGpaKNcKhcOXBJEoMUale
Zu4+4YoysB+yAv0iiPn1cnaHzmBaxDMmpSk5w3DkT1JGVne1ocJtDlOAsrupyrpl
MNenZVDmLMqmrXz+BRZgvyySCmbqn01Dh5yUybqhk2DXq8hFQvJrabUQMuR2NSLX
5G4Oq/wvb31ZT3MuWVBjk29Hp/8rC3r6Sp5aq52Racfixs2polZfUDfkI/rO4xU4
6s1wk1hoBoOolbI4xnwf4UFJRXuTOqzYS8UUJETUPTh96p95Tmd0OR9ywp2J3l+L
zmeBtV3M7BKEhU0KKq7LYXckmC5o+WGQzoV9s/y6J3D6ppXns6CmRnM6G4RQFIyE
DEI4M37S8gZEEWo1RQ2/aDnSkcfKbpSyj78v8cwwW57IShfH9OpmoXjwhBXMM2hN
qnVVTa03GDa/CQ8hi4MyvqOP/2EPHzLRXqQWHXDuJxxHBMeXK4Dm1YlXccCz1e/q
OR04Veo/GGde1EeqMrMcoxN1m0UiYDdALJrTl5fxxSlDx2o6dXzmTtbQfDV4N+PB
jlmSgll7/mBIHVi71/MykQdX5tljm/w11jqlt03saxKNLB68IhhjHnnUJsYFNZPy
fEoXeiLh6cOUjSCOW2Nc4A5zJcDO1QfHw2mUTy3V9ra+ta9dLJ4coiRqOglflw+S
EwRXrrBSdu4MAaJey6BK4GIZcHrTdtBATE7WwYLaNvQ9r5k2hYVc5QTcSdVMFKyj
TZ0sMwb0wakSCNINB7csRE5iDf2ATUJf1PsWRHXD9jbczlHbLXPdRy9WR/7ZAGwu
prHBPujmKKyrVCABi5Folw/Ag2fcqGEaK2DH8ftZ6xy04sPtpEIn2BzHbyaoaSIY
a88WOuE5iaZUj6GvYZoL9Nohw22QVrDmH7leixyRkLybesxKYpFyvz6WwDzoRZhX
JKdFrB7w1vOQZ/TDkQhwRijD9cu6Z1W2+muZjmRBnCuhRIgMEte62UkWVlOp/H3R
Haeo529pDzLkrwFVNZMMapjWyWXSM1hANde/MzBpdICGd9YP30nI0H+49hyZChUR
aX2BoXCXvj/NGMQu0K7fzNURpQOyF6S90kMpR0GG9s8ZvLETo6vToPsjAJdV2fDA
s4JQJLqBtg+SBEyRP8l/OkHH391AKzcybOScgubX7vJ1HRt4Mq4CZaRy1eua5jZ/
OVw+U2tKbJEkljop7AlJjw+23dvjpfhMjzS5LQIcPmF0oHYvE3SJEmA1EGlXh9bi
6aLjw5/9M8Qic3TpfdrJXstrGRS5eNlYRWD3Cj3i8WHej5kSSq3IHLimsLOln4kg
7LCYeFE91kxJgTWt7UrZ0P2F9A9p8qHPWElmqgLkDWG1KmGxHJ7f+RoZ1EGV4hag
fSzS7er6ev7GRTf4tMQRPNmO/DN1EWAWlm9AJmHOr8YJygsHPCv1sZZAh25Vy16o
U5DYpxmkwZ8G9rurDAmF1jUzYoyZoZo94b1nYu5jc5+U6n3bHT0e4bDQXYgCQHi9
g5AsE/30v30Tdk02noJbW4AiyPs4Rr0PXZs9ifyx3wCGdD1r38BYqDOh83C5Gqvz
zvRe5tx+Q0BHPxFGlJ3YL3z4sSgqZ0UavGVms/ck+TNb6AP8zcXz5zw7CuP7rZMq
89uEtEEeqtT+TL9CfiQdrpIHziLSfJ3TAbeIbmUWb45IcROM1OlYz1tN7R/NLcxK
6ztAOtgs/KR+eE308yQvDsN44zGlxr51GXrVG93Dn3jC1UFUVgIy53XeSD62n7Lq
zd79vXQ4FzFXp5J53crehH307JI2GmexeHJPSFuWdK6Iofoy5zmxoMBhP7W7nB64
uW4ImafFLzKY2e4FSjjkmNJUvDG27kJb57Cw3QvajBe8CMAbxlzjJQiLKFPxSSK8
fxWmkowe3L7jcEb6TTdHKqeLIRNICLI3VjItSaOGzqoQhtJv5253ImXy1w5xm103
NAtrD+WW1r/FCPX1/cxbfkG5VczKRnEdNtmcG5FGa+BRLagmFSe7v7hCTE9A235y
4SWwcynHn23WB3USASfy7aPmXLqkCjazcBGPYjbI+mnI/n/th/hU9qWvrfifpJTn
DzQ8kcggLRj1NbNogRFZ49TavkG7HgpA73YJUXhb5c8KLqFYcgxn0KK4Ym4yfeUy
braJxhSMzbAtzzEAlop8tiyGPxMt02RScL0XjRaSqap/ZzU+ditKvsnjbmEw/2Ig
unSQj3dyNYXvt0OqHwxp7U/AAKDzAF6SeOku4HdvS5ZI/+U4b3R+iewi0kt4NO/o
l9sF1Q6aeVDDa99FI7o4jIW2SMzOn00vSUKQ66rOurxYF0p+UzG05F0ZEAslsuYo
OXZxjH/aofgIx4SIMBBCx5DGM/S6d/1fyzmIn8ZbTnX3LTkTf2uHfOFpvRsvYZln
73cYRnlba3VpjKWa5EOVAL8pBUJ+XzbMt0sKpp9BdiN2S2XGPFK62wPqxO0KzMMq
eJK1YU6mSTq2gmDW1csh9B1Ma/0qvb/jwEEsh/G/Z2Vxoi+yDfj0JPPdCCQ/AwW0
6fD6uwq9/5ufINXUIuexK4iJmrWnAZ+waDXnQ87ugMyF4VizSo0O5CnGD4+jRN3O
o7glOKeiFQOh6QHnHDZ32hCHRWCO/aT4VGDPr9+byGf7Lda8rmOTNNI/TsgsHu9A
0uPwCGdmiCZPQQDDvkYWFqIKgsP3pw4+nZcB1FkW/cWODy0Tm+t7PpdqevOUDnCk
5tyR7wEsvzAxXb+kaHZ/S+gEMKYHEUFfutTxk1kuxyT4riwGvoMzKxKJKnfr7oTa
Dstup2khloQbZSv5LnyB5MwhgG6UTTH+yQkpYvmqrxQA2h/sbTiwiHMp321XPamq
eMSMPmXArhn2c6cUwwzTi1cgnI+yxLRS1lMSZXBMxvxKO+ogCCbyd1g4UOlNCNok
ONTDklwOqyhj8a+kaN6l8Aaw2SVzu+GP5pZW0ONP/UWQq05ZKKfJ4LeTeV/aG94F
fAFAZqo9DVDPU3HKQuvDgyfcLwTNhdmJcPEiev2esV41XeGt/7yJK4ZmwbaatiNA
V5f7hWU1S5W/k1WCA7Arf+iffzpTx0kmEhu1J1Y8tN7XflrWYOMZOxqzrsX5gvXg
2Rt9uNIbLHIGYkU0nDxVuZ9CHBvgIeF8sv/SAUDRXlUEQYSygDezhd1rOp0LCM+s
oIbzyj6AqRK+sqyPTidqAxtHG3ESxXKEB+J24SEMu1i6vRS1NzS8hJeRQ/trK+1D
x+zj6g2ap3E0kyEVNRF+RNTvc4fJUcYYpkDvk7f2BxbgknhFlKwkWTdTbcL0LdMu
9UkYfUVClrllrqFsCB9auRT2W0p2SxsvdPZOMDcMorBa5gf2K9Bt6635pRIjVbip
5TXveLe8OgfOFQPRg0vvnQJJ87nKDOmPcE1JznxC3fgVle4Bc9Cm4qXBcs3srtPU
PxsqgNrO46OziNTVrpLmcM2QOYfXtq99Qaz7JlrwJnZqZgDvfGJwtJxwCtJgMgoQ
QR0DN1Ifyz4XVtV05b1soDsqnY7tnPBpOELAaWQ+d5IFL/Z88kDN9VKVm6QFRtpw
UhiqSpzdDcz9llKcoeVrFi6NOrSOCATUepbk2fgCO0WN8pbxA35roqv3DiCJQheC
GMYwtQsf/s5ehJAS8Y5Om6s73HgNLK/syH9bn2SDO8i5LiToBVudzGtbXOIF5SXi
5gAZl+2qQBTOh5GgD3CBjeJhBya3+xzQ6Gsq1fNs3foIousQ198pS1skSc6XUdDj
qTuChGH+v0n0J0aocXEF7aemlG1fNEuPM0otIdKRUBYyw5JtnWOLL748HwjnEtMO
QWvzqbV9lIn9+Du6Fl1vz+nV8J+HCWSnE/75DjGrTLWnbA77iWtlAGGH/q9ven4H
y3tP78CENH1KSruKvufdg1/haletFMhAGobFRXPJqKRIvsfT+TDlWTHhlp0crLXH
DrQ087wRJ5vUYMSnUvX/k4UO8sxwOH4Sy0UXAZ+hY32J7q8/gBEq5p8b8FOoKify
h1JhftYAFclivt3/jy2QdWnjqhLhJ9mu8lxVdItN3TqxqNMFrFuH2dFhvkPGrbvn
cwXUzIuDsH8dKWI6K7yRrIircEaXV5RyGGimEqEufuLSQBk2slhbxCtZ5s3exdvi
VW14nJBvPfcEpOBPWo1/rkuL0t2varNzjqcQPcd4MIf1Kgmu5Q6/ZC7Qfqx4k/r0
d4A8P9G+Q39Aq0E/C8/GeCvoboJFYVC7a9JR9Qid84ZFh1Lc7YsPKicaV8o0wZlI
zlhwP+vQFqqYZlTyx4rZaBJjlf1EpnraRCkEQSjfTWfqAHcYRXvfGIOPOEquqhjr
hCKosHUkEJO2OFPWhUGQTucgnw5hCZKli3oDEUO2n8j83hyJBU7iKlLKinMYuk/i
dsrDPz9WQ0pD9IbZY+Uok3AcacKaEO5JGWumSMjF2QU7w1n3ouR9L6XxPCO/XPaw
yf+mRCkpADhaGYaPOlhcgp4/ZfDP6mzq81a3yfdjyKs0Nl/ubyy1ydiDdvUXV0uU
XO01MOBkOnrJV8+htRam4EEI1xcbGOiZTHqPkk/ZQXyozzEguVxAZI5QrVeiNsz/
fG6+R9c/vYKvotk6IBreZqhBleh6gau3Clk/5PDCSo+fVTxdgVto9H7k3KTPu2Uc
LqsErenYziJQZRCjNuCGjV6RIZZUSkmfCViPHACyc0hnwM+Y8EuPUkjqfNE1E89X
Ge6nQdgYcUpiCxSgSZ4wbqr20V70AX/RVoC3XsgiD6wxFHvMkdTQSzyEsx+T28sR
R0ELzUZizhwQwwm2iiZgUq73slwz6PbeUG6NkmnN1VEK/uK5YAguJJiJiWTveLSl
i/WnCrzI6iJ+QZj+WMGXnNtwqhyQn9myEpWYNq5YBuO0WSCeTEt9KjQafJg2V79i
TEEnkFDTNo00ek1qR8Q+SPx0EOH2WkPUf9SILeEfBSnQ4dvEb4IsWaG/rRN/TWLm
yaHu43ccp9AkV/JKDl3OlS2Wh2IZRND+er1B4srUubapUfTFl2ZpWszRCdZT3FL6
aCVKj1FV8xZVG7oKWFFGtHd4t6Ofq9zc4Qq00wP0JI3QWESqx/1klnBSuAPprWZ4
zFcqqyoIdGGvfDj9hilOm13s9G4/ZE2fThVMwD1xXMaLCqJ9XuCu9BYB7X34k7ja
Dqt8z+U9rR7H7k06SF+gk7KzjJmTuXPBYrn3vaF64g/WyWAyqn6J0u+zRxBbxZFj
5ptK+ZFy866uKjdhdZKR9o7/nHqYFT2S1ee8vftAKp0kG4ChCzW4GLB5LmAtCPZo
LZ2TSsBM58tSt2tQxCtUUmmcX0ocKbHz7K8yJ7g9LILaaAf8GHpzcOlpbfpvZdsM
CQ2UxfzfldFiHm2aUfLJkeWu6f10k+WbTobbUZ/jn0KPgBLiKW7LsxMQM1qIga4B
b7zsNcEvkPs56nM2VZzSDCKGyyGPBsac6SKryAteWLAbfjYlqjoubuAEd9Abwaku
OVN8fWky06F9rXYGU4PVeMgjwP6epS8AZvG4EY56DGbBTr8afI30xFbpZDmpv8IN
VnqVwnffHZ0dWL2AYv7yc9BTcdmBD+vhP5jg8GwRSQiioIJAolZX+sPPyxp0zbrE
wS4IyzRNBok8sMlDeGzA5Q2+YQNIN+NYxw1vuG6hZ03YJ2r6Yai3GUyj2WNzAnV3
kaNp1J8BPeSaRgAlEYo4HHPNGXzSSDd1pa4ZGe4jH9deVjN7inLQMRTuOxB7Yvo8
HPbHoZP4UwjpPX43TEMOACJxZ/hYJ4DDtHCLxYESuoaVmVa7xBc+FlIVMQR2/IX+
VMbgV97IJWsgIwmE2d+wubMwz6/0ubU36Xs56x+SqkUFdhk+w/F6/xmHLC0BZcUI
guzNsa9BGV2XDkcIm24Zv4m6Cx4Nm/I7AzotG/53OvM/yY3Nvr0bYh6trhGDNkuN
5fU6HBR730jXJGewMa2LuQ5xQnsQWDMgvfjTTQxkC5WqajilSSQ0onsEhUjKvxz5
CrN20FWzW5ZJYDoBugl9Oi2QOL7ZGviotEm/F7KmjOryRa8wLbzQrJXq0e6AZwDF
pPXwWI89jTSHlEu1L6wiCLJIjf1Thyw/mewpBhj+s8rVn4flThUFQv+IReYKtSXn
o12oCL8mYd7ReEf6sZ7DYpJgfI7Dr6On+uSqfMGlWUV1U6kmA3qPqBRulyEbuXvg
JaAENyBfL0zsFE2KQ7upFCnY3oRe334tj4QVHWMClll1WwurVM7wx9njpCnwWIBD
GT5MOpfvm2e7jhEybvsU8ExcWsW5tQ9P+WkGVewsLFaS6hKj+kqNLWQFNarqfUfo
iSU1c2yd8wh8wAH9gcxzSR1NhgUQ/wSikaep56QjtvkecseZQotrP2z3UW5l5FbS
voruOdTVa5wykssHS4vcu/Wx/YzY6nkFkSANLjSG/eVks16oV5e0lzqg1SH+zm9f
Ap/eUOoaOqFI/wDWWBfmvRPO07O/NrhTs3kKFxO4t9mpVHPTx3eH7ZoY3C5g+xWF
4ETj/+AnBvRgFH0MuRHPmkQnXDFKhJUMLOXYRYdani1NMybOlbEgKB+AdUOshqwW
YP6c/6pArE1A+dmv/cgTz7PSlioxgQeuTXcaW/TDZowUt+8hXFX+PA0NL0BkFP0d
IPUxEtqT9XY3wQiElNrl2Xyht7IwVhGqQ5ieRjHFl1LxJMxs4PR3CwFV6TK1Cj6x
K2h2SeLQv8ZQ2w/+aHIWafeM6UoM/7aCd2+goCwtZkWe2yHHsdVZXZaYpPEoxl1Q
A+yUyKyulCM2W/fLzXTJzvrPy7zKA8Nw/rn9M8kvp6R2ZzqcrvrfO5jOD4FZu2CV
8bN4/yGHe3BEXl9P3tbgkHBotOXw6EOrcRtpdmpcRfLTBWw5EutrGBNtyiYpL1xo
j8Z/BaizejSFidRJ44mXb0WD2QuivfIgoDvOEDx7dghUXN228I0I5v81lyZQZTFv
+RP99qXLxOb9LYnvmLhb82bLDEFKc5McxPNzjm2I83p0VYBNOaquWPOrxo6E9xji
p90k4ZI1s/TDRQchh1MqyZIqy3WIn7X6wfs+Eb2BzLG0wIoDAry9PEcBQSKLj3N9
RuCNIwM6JlFVNdz/lOaCUG15H+97yUEC/Cfv9337Bfkr+QOpfic3hFF913B/AW8H
NruY31U33juH9dylmfUul6LkJUmQtlyG0RWfqap3JZ41/jdQBLwjYfsWiPZIDmY5
UILiJ8TmLuVOy5GwPuamNYn9POVf/qac7QEfbwv7vgIfCguxJHSXohrb2xcbf62V
lXxPqnQspplAD5egtyHfWvu6LqC0TbSbdlyyGDt0ofbYKBHzFiyKUHfggkY/VhE3
EfK5TfUi0zqRele7C6Mokl5X0obAS3mAn7y9t/0h9N5NoOZpXXXoYc1tBy/OL6oP
O5tXt5HFMmTb61i3CJc8deYBU5ZkrR9KbAgKC5/23yx99MqoJuReuqK0ECfNQnhX
ORO/M0pzkkXNVXpFxrnojE8qfNKJyzVYJpbzW/YNJFZov7fqm0i8IfWPduh4H+wh
2qutL41hJbM7fkF1kw918+abfHXz2UbOwJEw8JaHgxU6wHDoYygp6X+EBcSubjPK
GxdlhAuWBHxXHN2as2flABI8VompjEhmAwMUHJzz650GLIm06GYTw0tDa4T6o+gP
WTBKJ1QX0Q/Zq1zSJZ6Yamix9zJxWYDctfJCvnjPEuBKO4afmMy0c4IBMucZJeDP
npDXcUev87vlWk5CcJ4bxM3SxgptjgUd6A0MS9Nb24qJDFjyTOM3pSfry/5E4IOG
P7fpOeiT6a7rqDtzvhuSi+d1HfLPnmGqw9Fi79VshvBnZwTC4BMOKI6FLTEfwEHz
aQUbazEgB0oAn1DhtEHEOyBDI9biW2eaPja/J7hv3kc9TW9rqrpFaWrRaNVjU4Xu
jLEM37P/wNlwJ2wUP+4OmMVMdCshj6NmV9TNEHwpwqxGOFqVS2wlN4n/Lwmwefmz
NDnWMaYkWcGrIf75sfvBuwSyF/PBdmMitibRVgDAruB/IvBZCQtU/SE9TF4/Y7s4
ZOsxOE0mIM2G+2qQ+CnpnS4LXpvx/lgqonzp7zVFgtg6gvVa+Nl9FAO86MVu4Lhl
sUqVlCDw9mxwhyKzICU16fgPsnx43+HLu0aDWGJRNapto7pO5xTyXZv+sk72GNwa
BgpOzrUR/gFW/b+PgRnSE4uT71WepIixKA8qvMZ2VhJ9/EUgF2uCd7xVXMn+L+cR
HuB5hviIyrTDcddd/bUjpsZ1JDuPw+mhO89oGNdPbFrCGSQ96YnACGm58IYnRsit
fGj2M8Cm+0SSWt1a4rrXc4H1PiG778eooO3581wFfh3xeToATdlCjCvXPatf4RF+
qtdQ+QbaqWSgvYGHHSKxEsaH0Yd5DyzS/Qp9ecMYP9A50rkLfRaT0wZ2lxzHUrxW
q7jSSpOdbWRzPVcVDFoEbnpfV0gWNotMxLarJlEGVPwVhPRGjDfpLm3dTkNzy2cP
m1NXKh1EETiuvF/jEzHeb7BzydRU+2t/QKpDK4+bZFfSuBeBJa+fYOrE+s3rqa00
2etfp+RimbmLVCDZyxfJu3+JYvP6dFhPlfp6blUaUf2gD6+UmnhpYmZaazkPShYe
r2EiXvfkbJAIpOf4oBs37iHj0fko+ArFY1nvrNkbfMUJgUkZgoMLeWV0z6IUXfis
zCGw6b/CYj+zmiEPY0Ji7jIdT4kb/gQWJ3yQj+QcpKMY5xQqjU3GVV/r8RJoDI65
eMk7ovU0tm2zoCT3rjRCUzo1cwrNbihQLVSqpNPBF/ZCPZPWKRrQawUEOSjMvOm/
oW02Bql9UsNypT9uoHxalqHIUIij5JNtR/wiQUV93jn1+FqdDAlL8GIpkMtBxQda
vzD3uin/qoigPmyPPc5FkREKSolYa9QDlpbBzjpa5JlE4KM8eVoTw27cMTP9T8sP
aIrSfI7DJji5dLlTVVmVKwFjLCfe7LNcYh8eLOe1gisX/HWrkohfxk6vWxkgZrIu
Yi+/cDwQXgtx24YumTYtsISYjT07zP2Pf50JbmG6N2nIjEfQNJWWUjtbAvLBe6MW
VuOs0WNy1vOI20a+SNmi1ToGtPGgCxkVWO+TlI/2U2jLKREmas956RVhstdncGXh
r6bCL7mv26fBH2mRgJFF2MOBab9/VQCE8ZTPi53du+7vAUwUmsALhLT1hheyFimy
2ItDt+O/LyNu/xadml6a7oPtFzUQzyRaQuUyT2oIMGgW/C04bJGEWKCeqd8Ars1a
NupMgCrs1msKEuLHdlHZJ2g9IRPIAeoPBQ08fP2Anzxwq/6tFWDE4ipjJ4d3igBc
apZCH154EfSQAc+zNPBtoBv/SO2FEveFMrlComcnLhk4mbcOXkIsopcwCssJBeE0
lCAp3q5pKEfLpV7UE2i9HHLPKbkSW+1J5l1WkqaixQFBQFOLR4XTakNe4yhO3cPC
VjNzBR4PEkNzaRfZ5q4bvVZ39P0Iduv0IbAIVBRY00EQvE8xKENKhiyDc/NTL5vx
smWRYh4wvhGsaYmkRzIPYufRSXJ8dAxiD80fe7LJ9ttaPQ+R3GN3RmvSmLwcLbW2
vJfUB02iF/S9twd217dfRhW8tQFMa8h15B+CK/YPdzcOHm3LA3PSWVgFcFgwsM+B
A4wlnJKFM39zsdzm96k+ecBlTg/JGWgNBRQ7V+Be11CMhG3BRYGW6cD2AyfCtZ7o
kT92rtOSgU8EYNnzDcKQBCorxVoaIU4/th34elKVGd4QSHbSqNJtuFzuQ+0uipVY
/IoQFAEOGGFet1OsQl5OAXW500X1TJPNeIRbD4eXZ7UH02hO/zlxOujthp3PNEA+
xW6DClcxz+6CiQmjQVidLdRFjpNqlzRt+rRbL8vcCx5gB+iUxD1sFI7kO+4Qs08I
se3Cq3MvRIjJ6WfJJiVNOPr5F2G6V0QQdYjq9bv3wEHNCEnGXYUl1HDMabZJPhfa
u/2QbSkqgEiaSvA7rpUEhhLg1mIopMg3FfbyryKIutbR7c12RUoi2cAkBssWQXC8
5Kx6WcXjXGlc6PHZlVIPOHDuVl/zuOQxvtGy/vynPYbwE5Qt+ZhyGf4H/tbNZ3Zs
uGCzlomy0NlUtm6NdNTNWUyPD0vdhi7GYNwB9Crwd7EdY2GwHC5n0/0BEDtxyE7E
VOcWRn+UBP82Hyy1jwfDA6Hs4pEs5n1rlmK36R3SyY0/v/+n3fuDA/PoFoXFdrvI
UfLIcD+hsX8GGiW3/dqbxXTiR49YBL+CEH0vKuWulQ7RqYirT3FYauPCQgKE8spt
+w45yHCWf6U48ijg8qR+lYAcPLrfxChn7CRLn/gJkXMEW8FHD6fSyKehi+pC2MvY
n6jWTACYxfhMXOlcKWBxGvU1Q3lVDIXV6HPt7t+km6XAqz2MVYPTpjPIyQndFdpy
krcWtfRdX/sTG4/IKBCK4+WfNfoHIygkfHxB3JmY76Ism1b2z6oY+tJLTop1cYP7
3Y0Lack7AaNTu/c3bKqYgNLsKfT95v6sAMWS2Rx0Pe6Xyos5yqDwX4Zm0FWOMhfq
mqgE6wd/X9VHLgntbrB8SqSeOr4k0gRIHDf7OsH5PqXwMaLGJqeaD3DI+Jx57t+O
SdTkbr6NhVWE7970xycR0WyWNsDsUSEOh2/JaAD12H5NG/CnWLHZHiYFDOMqA/mI
8+q43Y7jtJ9ZZgexYTbgFZ0Se0biYb4f/2f8viSkMrI4DxSrV4Co4dRdJhMgKEfG
6N1pO12oDU1wxGqngOS2v0dsH+7x9c32JzkT5loMeWVJzWoq84gd6GfxWqWUNJOb
UHjpAKPx2BGhrXCCp4Xln4zwBG8NNM8tEnUPO8dzaDccvfJLP5/xir7iD3kD81zr
4xwam/dm14j1rWzXwTM/N15jwGGpf1R2U+5bgO/yoPvMh2F/6lCjZyOd7Catat5p
JRAh2F83bDOCpBJJERLcirb3+Uacj2QjAFRGt3SIMS7AFZ9DKCsbkGSU/xwisY6O
ICMmyYMpDTjfSRKrelBPeMfJSCYf3G4zV57Ta+ZY6IfvNwHmsgFcXhHc6wpR5ulf
QlEUvxSzEtJ385Df0X3C9gEsmFuMSn0V3K9Hu9+k2g3Z5AvXUg2qTGtqD80+G1dU
b0SLy7NjHoCtQVqAsjZMMsCKQSQgDyRuH/fKBia9r+22/1ZAk/M+MsN7C1clBN3O
d3dqDox8Bfide5zVr8Q0d+Oa4jEO65g0QwCQMP6B6zUkx/UI5YHJLc4/DlkIH9I4
fCY3O/IDSryeHeNdWk3Eg1yx6nHX164PU+nc5e4ur92OcjoR/EoThk5f7FxServ4
LUa65ScneFiWBmNukWgCYmsU3EiVenIFJYZEzf/X6/KLI/w8BIpfSiPHh1dH9gtq
OZJwX2oBSa1kAltuePlpN/D+GiaT6ZjkxlHzr9YYFhSvT/FvVKzB0fG2bA7Mejq/
p5q6acA9ESHcktCYzusmJg/xeAaws91l4TWHApkdkl+kGh4vYuobBsFEqkSl3LLG
4amsHHL4lK7rbeIuPshDSm2eB/V3+lTPf8XyXCfYa8DEXXt8XamXql1a654a4qCS
CxXxB1NOpsDyrX7AWa5w3IPNln8Jpgi1MiTq9F4PBOPvVhjT2Hs2gx/AmtQurlEJ
dBPXFU3Hw3b/6zmJXPT9ooDg2OSLgcliBtlpa4rLtRK8LmtmXqnomF1fLKzA9Prb
78fadFBJF33+0TjeUTMvRCWC8BYuuFHryDygMWKAhdswh1+sRuM4hreFojayBF3k
jzrrwC9NtbVCCR2zoLGeQCj9yw6y0q/sbZ/qPENh9ZcwJFA1RdUc1b9+mn+CWom+
vdoUADKJscnuu/wP4oXuKB1LaWphZXGTEWaDTQk/C7D4mKWwH1Yc5h/ZZMvasUIw
FYTmN+UepijWr+lpaz7XHcpE5o4gexyRPz8R6SgdYhTcNscMZ7S2gWRgcfJ9ddjv
5P2HGHldG7JTQpNyH1oYWcWB5lcw4DF4ZRVr2nr5E76BOX/13d+I4X7gqcloRKgf
tGav3gdMSb6jDbQYONDXIMPNRJdyX7PRbnWwYyoRh71MsukVjSHcEYHmTKGCLZXm
cKLdEyVO7VdQ1/NbNNXf8OB/xkL/uph7iK5MAeGBQpbZjtYlWFWlDdyB4CAGZXc1
qKgiED1NQ99NX5Wz2ZzUEtkfWJDXispu7IU5WPWKKPe8KOXVSTK/gcbvHNNhl2WS
zVpF0Vt51wRzqu9FB+gqD7yw+8SJICMmwRKHwNNXVFojPZPIwAZ6RHnDWbz5QqtV
7bNUQIkiuRAch8yU6g+aSGBbZ70R3iJeGcXAL8N3KKxEJXnPn+7FV0HzlF7027QO
eimdUDu1PYe6RqkLblQkRYg8dkSqMAa+jroikIfBrK7RY/1L0PPIU1YPOzlsc9At
HvbzVSnJEXK5SFb4kXsl8sUlRL/qWBcmRnopeK3gfimVfSb5RFGCrFScWNizbfuD
YW+jzi8Opy1kl2299/XieGoRHA9S4Ahwa3HtpAlU1aSvd79sBv+nS56PTKO9t1ZC
Ndvdejaedl8+jr5L3zwahaFTqJi2/MpL5ISOBkZILxe0T+f0lcyrNjmE20ct8mJ8
HxusyCs3i6RB/P2d/x5WUQ/MyBCGTVyonmBrSHoracgssfFfXXq0jec7ICXLuxil
bSEE3Kgt7auXEULvzSIgfV+ZOkH5z7vmv8mfGtOI549oRWhKnYuK2dahnf4xr6eW
7yLx4pUEEPMa4GTzpovui6At34cMJEhht+uPZXNkqLcJrb+LxmgYYV5VVWC8uVyF
UAXpQ4lxLa0NYRDoJLV4uLIsvs4ioFg9tnSW9R02TrUK/xKipb4pcDwMyKgqKBn0
ItnYRk/lIU8Rxqhg+3Y1kUUj3AJMG8xfHxP1kz2ktMMpHoPxbKHLGJzgXHVtFZkG
/jMHobw9OAOZQBdRwLPzUMBLQJAZZk8O1l7opt0ZYUPqtISEdtK31t8xlAJ24uGy
k/3o7JM1t/E5QKQSCpOcl3hn1H7RoilIyWb5llBdsC64abAEp3/mB2ptNZ1Q576c
Jh8WaveZIgeSIWF37wwdRcnlWJjJ22ItKtWzgLdNl9QOorl3eGL5fmV7oQk/w0kV
wb3MRp6+XFfH2Q+nLMf7jyBt7WBNq2yASKx9hkiVE8stOVAhEpRJlHflsdVGugxF
qUr5kHcUQ5UgzFBJxplV+kIY4KxgclbJvGU3QjZo7qX9xmzoncSH0JGDu5XnsWPN
PqxK6pCyWa+uZxTb/A9YfVUPyJYdwy1fRxdUlCm2asFpNSEgVKvk2WkielLl1IqW
ug5UbQ5zlCQfHikO93Uz06iHA0ynMZtBZBCihPdVNp94D3v5ELOy8rVp1l9mnNoT
vN3bhBJBkdZlvCcrg+GxWN+q+DE3ZyBkPxy2dTt9mcvd0ePewnlmwoiUwfa/dd+d
ipmJB6DqlpMECByFEikSuB0uIxT+KqTuExfPVVbJTDdnUAmNchMpz6Uj/hhnVBXz
nX8BzonMG8KtPsh9WhOHL+3FfcuzSCSCjCMD8ZDbZD2C4s1LRLD3kr6vLj/HfeF7
t82gC56D6AIeKUNK1vXx9MxT4C9Hz8g9NA1K7BBvjDQ9bU6qhgqskCnlrj2VzoF2
2dxTrq/RLkbvIhaOoXqvuSyoitIyyx8G58l35EGVaFK0w0cMNrSD8vYGX6h3ICEi
1DJU03AqjNX2lSa5FNCr3hmvTNwcFOvv3I/7jEvbmUuL3cr7xoApedhPNQie2I+c
Ph4sbwJaTq7l9LyEN0qI9FYRAHkIxxv0wKcuSogcGCMnr/pikno6rQRiuZn2Q/zq
tlh7+eWwgh8FBhziCtwqK93SaibzLQ2l+dyKyZf1xwbXTLa3IG6TKJbp/+VgiwCC
5VjWOl0Cov1t05nuoFJiONXMc2VU4SXEhWYfVH49g1eByO1bFxC1VACa2cdpMggD
J5Wu8Ts3C2sVBRYcxMZkgiQUYTHYjnMrtVH/KJww8g9WqnevxYuAKk56XAKXDqQv
Gk5JgYQJ9qgQSpZennTMCkEQVn2ows1kwtPEPTz96tXQWtRbwq19F1LSXPqNcCNq
WFA764Hw9mS7DoNVwtnxwYn+hyX7Fj3sD+LKROX8kVK9UJ37QkNdlS+RXDgxE6in
axbJCHxC/gL6NmpN0P+wM6j5UQzAGjIsc8JLEYwwq+CKVAK0cAXIE10WehmdwHor
ltfdu+T5rSWKoe6XS2klBASwxHuQMGyU7lNYExnFgFmB2CB1FbaKo37SMy62Wmx6
R/xIJMpEP5uG4Nb+kIFzfm0ent5Sx3AO6GEWfOxAnNuDAmnATVVcx31wl4IXTUvA
fCPZWkjbj8oCZi1vpTWibEsI8KS0Df9DQmSRvVwjBAm2vdfyzPb5M0hy/9/n20gC
Vda6ZR+SuCoUzKQGBEM+OwcnbE5ZbJVCrk8F5Lx0ZhIw2gsSmKfSMZP/68xZCYdF
GQrLbUv4DoOQVU8YOX4pLYYiO4rWoP6xXApBvFL0rXoWGZAnsUCo9/9e5AB45i6q
TdhnqMyZlwxXI+EsC2lv4U4IJpBZjcyquvvQPgc5SYBQEfGoS68faOxWjZZaUjXA
K2KJTjvJZHdZ5+D/e51F+soGER49G7EEnDztv/py9swKMD0hP4DoCJEbURu5WuvD
MXj1/S1+4vGVSMfFfRQd1JcRaDKghvU2NjbUguv5hl88y1pqgyOaWxslyR+ZhiRa
e18VClE2MUkcezraNhnnLizl9k9ev9CQIHfA39zCseb0WjTYbU+9+7+GRKloDU23
DLcOSf4+pmj3XpWw0xwXzLg26DXsIqJc9/SfN11kXq9csjjjO7EqxfwpM6eDqBIl
qcZ32vvSpX0tqh2GJ1L9hdqxroqUP5gF6LHHihV1hJKmW7Stg8AwI1035JqSuEKm
kdiYtOO8iHs4BHoQ3YXNGlrXAIMXLm5Q33Eb31cKRHLxyrm7ShTYLm2wEqbkN1u9
cJrkMBnKnBpZOAw8YqYLKmrz0+jWqYaASxTaRskyGyOXBMEhT6Qdlys0F8Z3B9xN
DUy/gpGAy5F2g2abjmnIHXXUS0ZEul8kOCYuTmJwh2r9RRsoThyQu2RC6k9CKMsA
yZ5+OjXyj98M2ngDV+xy7DqWwxXTbVMpTjk3y8cBtoXhMXPAUKs2TFH3paKC7Xsr
r8AgESL6o2IMhUWviwo3UiuZRzGmlRrNAYnzbQyVKx371XLg+j3hP/Jleukt8TKI
aBh+n7m8DDKJTS3ubaLB/EJeSa+EBzGksITt2KrmBLaA/sPVKVBJGBUSGoBEnoMx
urJpj/v3qkb+Dulkb1lBMyucp/B7ZbQGSba4aY2zybMOK9EEz7pN0CVJ5tunojeD
jtp+mZsH5SmHPKyO7jzcGDGg527dKkl1tbh5La7xUdvSfAuQj3WpzDB5YVjd8Trp
R9IRg8gSGKuApvx5SHSvgo5+8ct8dzTA5c7fZoWl5mB8bMZbkbS37dLtCMglhxrQ
OLqoQJNEmRHuDlDCHQ7sR3OD5TEbgv1IVWRmxYv+C7iR8f+/IoOe9d4uKo9A15o3
PtG4EZXSUS8EAE5U9mfs58OFV7tF48U3cHFjdfiMVnAy3DCp/+oU/ZphHvAdf4Ye
4hA/7nDAAK1kWH+XjhjBhB/qwkqs+tmWEs05W4rZOkey0xid2tgJhTV7D8ltRNb9
t2Pbjv808Iynq1N19aG5tT+Htn3/JctoJH/wIAt0Am9qgxtDHC6/5Mh7jaZFnVSM
oagV07tgqkULuvcvgvidWdcZvfsnCcVDqUkXEtkE7PEOnVnPX2hbAdjVS2iEddCE
pUY5KHuYi634PD4i6/Q1TtLqTWBkYq6+2MVkipybAgRm51eSDjPFvnPBVOdtm9DZ
itidQDAJGmohAKIRT2o5yhsTvzDgtrM0JvuF37ETaCWLNJbylV/ezqTKy05K++rR
Y7QPZaCNrd5HUoEYXWb8MMJUDUHaI353+DSDHddbVFn9zKSjsgBniD2rEJpw0CVU
dqClfDcGB6hv79gQBb27c19Q1MdioKmnwaemXWDj0ZkMyBPTRuFz3+IdN3X2T1q8
gYh7WQYlo7VTmbSKFg/EVOKHgKxcU10bKMWNVu3HQWXeAqK4u1V0Qe4nVjAojFj0
fd9pK6oEwl7b2j5aDk2MWpPVHcJfeNtJHus7xXF8vo53OTMBjxZbZqMaUG+99ijG
pifLuYRsvYH0XSTm+2LifExJmo9LGLVU9cOWhku82QsN9LbQxVsHePgU7WQdPRQG
wzczSPQG1/4B6FLHgjDwcM2ntg2Kfn0Yj15HX2lQevCrattIcRYNtQaOF7vVLnTw
cgO3+4IqIfOMsn72oR3V9y6DDeSTAY2d8e60+POh6xwrTNq3yG3q3xXQStkpTlj2
w2h4zXoY7AgAGiqKUG7TYEQ27jgVGPHXopwYGERk6JnfLRsAA0ErDPbewVuh4dfn
yLVh4A9ICFd6ijSZ4xf5TgAirotNtKomRGpRL5rCcWYKBYkRcYhMWTmzG4iKF3au
pIndCel5sI17lQVzYQrVqmUbXolemtPiTWPXTkth7wBo6Pqg7yWlQZvjKKfHPStW
kpUMKantezEqDZwzg75IEKErnc5weuEdqmiwNKvR7y4Ya4DR+kwpMV/BQ3aw0+ag
3xYZBDV+AATimZqUkSlknloeSWbDL5wCWATi7+opr4KixzV0UIZcDxmPtcBk24np
YQSj8f7bWifD5wlesjZUIBRc/3wsbs/kuEV8/UOkw9QE2KsE0y+oDMKbYIJRF7Lg
1l27NyFP7JvpxtP9F8tkjHMLQu87Q+otFW7HmTgcnRFZ0jSGDCnn+tqTPWc4/DiS
q3B/+IwDmgRkBlDaxrLs8juOhtokRXb5aUcs2OvXy3HMPYx/2j5ou+Uh1dxhqy06
ic4kRkQOOc8t4oT7KBwI/hDihXYr06JXCiQTUnagGMQLmOrYdWX7seFVMdPSXm5b
yEOEH7k8RJYNyBamuNOlMtuOAm8PxH+ZAK6Oi/BrZFhMXuWmtqb4X/xp+VwP31YE
29qKd76Y5nrNjIGtqjt4xBIuZWsvjKdWltU4nTD/uvmqnm3bP1Mu6sUMgY76wkYV
pJUDTFytgPchp+1wn8Dea+y14Ka8FOY7ztQZv6wCNStV0fVrxRZQ9slal0DSK4rK
98b62GVtbmXgcLji01z9WOKXvi8bKRMBSRxYlCkmCVnrv7W535FNiDfsNT5FjmT6
ie5GIaOt8UVq2WgWVcJszfrQGqDoLBsATpRggbO677kcCSmKA5iFIZgHdI+2ue8s
pFVRhTvwyni2PC9w/NhDvzHImwRxV0vzH9fWgWEUB7rOPDfCuvooCSOhW6KozzY8
KNXJ9w5sOan6+lO6b9sfJZaWWLxXNlSPLF9tqb2jKUdI74mFQ/RIWf0JG4YWE0DV
d+RJ8SOT1baHGNS+M6fGLBudmT7odHfS9rdo0rfLrxvx47ICEpVuNYnQkIESaRaY
yrSY1Lzs/vCH4ZqD6LHT0LNbX+m2c+LQSbdzqYoq5Wd0Sr+zGxJOVFn5ytMp0N1q
1ZWwXnqnNkGjqTd8gxd2W4PD+LDNOHg60ph4A8D+rpnO/FHs+6VHfLVw8XQ7O706
UIFpaYZDuabFJccBvuoC7w0wPh7mSbQsjY26hnWyU84b8w0Qc+pAIz/2lgc/PGTv
0HmDVZm1AnbZ0TYAZEteplFhRdc19IiGOklggzoFlgGKW0fDX5kigy89jlhAUTKK
EYyZtbb3G6QXdfkYKVuTO8bZ/jrycnyShNgKT+tznoAx4Mu1fJZO6kzFoue/qFyd
L9yuZOpetSJ+zRsyWjXbmv4hodN2SYeuqszG8T6xcEPr53jKuAZhSnGkOXrfUpjE
UrFB7sFu5QHrdbUJ4acNCjCPI/CagPvY8fysc+zbjmhpG0NKVnpMGD6Kz+CfusPm
cMun/+7ClKpIg8ZzJURqvHeikJqpln/cCMbTEWquCT8JyiUihD4jRCTq6rIf3tVt
s0wUIk5dVkwB/SA8tHX0ZXKrR4FeaIzPpeizERVmWtL4beNfY2uui+ESq1Mb1bL9
K96w5iM92ga8olhOOUvW1vB6S8IE+IlFg4nOYL5SaD4PF9FSC/kJ9O/lUfJzCkot
d1fS9G+M1ThN6OAOYQKrvPa2nh8tiLC7MVz1i9OwRMBcJCRMJ7r6177Rs9XUK69H
n47RIAt6MH/AM5ebtxG7aO9RyVlyjroba2YvFc62pyQjkCdibxpTSG5pzMH1Rbus
O5hBilkDCl8G7HgunjC9uOQ4wiwdrr/wEITdu8vKcIZPYSaA9fVsk4KvLfqCa0am
MEATGReTECGnJwgwx6gbDEYI9o+ZG/iZraMOS6oTCZDlwt6miOIWI48428jdCNnn
TBc4Rb2RFliFmP2Z9r5eX6XF0fla1zwYAU5d2jKRTTKnqQNSjmRySKOwll1Qq1rg
VtuDkqd7RaGR0LlrEU1bPH5H6VEQ7YPTcNQ8yYWxTvg04eXT71MT8JdBEt6IY4OH
BGnczW+6l0t7kw3/JjI0H8A2lL/Dki8lT7Ioff1r3/wShnCHwrHVVyR5yYif0NpD
LbJA1YiuRZwhwWU2fTClm3B2QXS2hMBrRfcB8uWf9/onh+6kMwe8CujgOVOwGaT2
K3bqT84MoGtuvmyBVQmynj8JjCIZG8zqO8yYJmq9Eqti0qVkg+uzV0L9QSJTG+uJ
ea71uW9X7f1TwWU711dWa+2dTUKoTDPayOeXqCdqUIRn5lFks5DABbkQxJFr9c7t
kO3uG9Uup2MKnBc76BqIAaiBj/3Zfiv6f/hsNsUZ8YFoAy5LCqO7c9mB7YxlvF/A
o3ULbtefjU977mO5/jomDqst32UPAKGTOGVlhCYMli8Jxen50mSUkTWkhmGbKnjy
uKGrFacQIjnnozu/YC993yvh93xTku8AfULi9AVQprF/65rtm9JFUjVdTmElX5ys
LXpeE+JEeu6ZF5B56HcVaXXAzw7+UL9g+6DMmlpX0RQloZEEdPF962ssmiqY2ab/
0UZ0GIk3V4445IXxJn1t3v+3O+uX9oKeXFt7RjQN+zT0x90R+gX2TbcCm0UAJOVm
uNhIB9nR5GlQNCvMCEmj4ixxVriT3+CUak7Y9wAJv5CJYi3NaVgvFVHpOZsdB0do
LDBRGdleU5etVNMEIgnuG1xJWrx8sGC+5p5a3ufUIvLhMQ5UFVHo8/sAT4Qbylj+
3ajBVon9YvT6W9ht5AWB34aC82dd2KmdCV4tr7nJKmNXcwG6YhX/8DIW27DQc1BA
Jk8vSTSXTGoWdXibqoRYDjaIUjBnAMZtO4RpI2piAD9D9fEfNgs2cnUi6QaULJzO
N7kbg+AvUsZ76pQGSaHaFULtnv3v3dkV+ALdIfvP8MoLjKQjoMT7D+AZdOjIupl6
TQo12TzEWWhySI+LwrTBeEc3ONEUciBv/0Ir7y4AboFn5k0DRK1/0lUZA/J+Vxfv
AxNWogKEYqNHt1vZTM+xLvMtPM+cKHfCHCNnCzTeNirNv+20GDdiFIKGJ3jldZ5s
+BSdI5je9QZbdru0PFbPsrtU45bnjeJOaoKXukTzn7FqbZKDE/5wm1skWoPNHXMZ
skmxfOjA7VSiEo/GqxCty8oSr4oimc5+EcCVNX0tW2368+1+QZEmSvLyaVNVXJlB
PMUEKcUnh0ayG4ncKPQXiHtDc5rKn9eLV6avOrgFESyGqd3QwLcj3VTb9UUzgOaS
8RHHHiqkaS+7ItdpfM0SYWveaV5j5x5tA8VqzhBKA5CTnQ0W+bt07YF908OeMrrl
bsYTQOqab1ro2dOuUqf2qw3iMRY+OuoW4bNZWgBe4IcXpQI+r+5Et0VtvZvoEvv0
BCD2XiFVNaKHV1tWjyCXG6390f5wN2vTqHp5PDdWNAo9n3Qm+ihfTtn9r/k2Nagj
AMfnTl623jJQagM0ynUPQn/rJ9YhE4udTm/BL2BdAMLVoGjbgc5PtU226HcQLmy4
uSiUQBpeffdD1ayJAA08BiR/Zrj34vyXi8P3CZXrmnfuiQhW3JkyYS7OpVWFHKiH
AoTpIHhm4604gRrSHec+z/DwvVYj1ct6Il7r8Klg+lsGK27bt3vVk4k4qwFYmGfk
NzqEMxwB346Iycc1LDXbEkbMHZZVRsDg9tH9K4jXVRHg8ygElTbN8hQJDazsLRHJ
pqatvOuyl8YMoBi8D9n1VdUpUyHrg+dRzaJ8pgYPPmErpOVwJP7RRO6+OSnVBUMp
1wEIcGcdrTKCKiU/guYUs92IfLUTzAK4ZHjICvOTdosPWcWyTx8XVetKuJ/Z3bDa
C8YgGCrANhM/6phiupi/vMY5y3fOC4eZ+fLIO9fbbchv4Mfgq7zbIBCF4/fTv6/i
f7ApIcnejerbaliOG5RPNWwPztEMdFl4+zT8SW+rbEO20/RZc03XC3lnuzKJQzRX
n7hditQU87Y2Zv1pZOol/OL1CYodQLEgEskXI6nZ4ZkM0w+pdYaLn11FoAcsmjcJ
yejR38MfwzvmeG2482UoET3KqXV92AILcAch09O+Oz89F+JHeipZ0bAsHLRVC8rJ
e7nKUdbZo9OnjxPpvlFEP5ZbcsjXKhcD4/+G8tuQ4Z6ONGRb8BdsgPS1Iq6b9c/w
fh3kWbM3McVgGTG4BzBerKu+QLMvtN8PKji6PdefHMn/rDpomvRMe9f9MdxEy5TF
lZXH/lqYA947FmDC5410Yt5zYwmSR4jkal+YKraD4ymJZkhPnAeiF9qRgVV7XiUX
wrSgdRDSWRuYOznaQC40RsJyjvCHBr1jBGOk5YA7DYRSm1LNXdLvwTAJcn17AEx4
g86rhaKSveRbGQgE0/wrfdJ4JddXzowO5qsZfgPgl7xb5JzjpDl2Aj2P9aUVS7gD
I+N+Lnnz7m7FzeuFvXBIDSt3B5bI/Bj9cfPNd+krHiqXaFfHuOiYpXN+quViFeKP
mxvFp5jCdCaLi/cLg2Oj0Fm/yrWJQYc0NplSnuPScJIyJPP5OTsXFn43qWChZ5Z8
y+ojCHNY3P4ZkYo1FFBFsIYvye6PCkc3I5Ws9qUdsxrd7ZcU/r/RZ6YfyhlYDrDY
0/PqUHUD4dDcfEQzmvhtE3J5D5vO5FW7lCJm2Qt+SNfkPz0ASa8kG9H3QSRXm7t5
hhv3G93V0GJG6Uqd7f57PhTKCinoLxE+FaJn6qkQcED2ea01xtqDSaCshhWsPnKG
kHpjHunn/AFlnL9tWMQjBHmr4N8qeZ2deWJnXGMWT6XHqSBx4cjHi1YiZp+flZ4c
YmAy7Z9WQhdbzwmt9W8N9Mqy1HOOeSr8WWueAbtOe7P2yHDvXO6hUrvf0rf998VH
EnfcnzDGSWWU/kn1NcYpDBD4eRDTpzeaIEJapIjlNRhRvTsglqVxHv5NewNvINwa
X8iscDD3kaHV3stMwLkO+ZtI1PXCU3uZR7uQ0GLdq4pCGvm0X4g8eRrX/ORhn4Yt
YhqfMSxOTNWlYMIvjo+zgjeqUO0s7gQjNVog9YaCUBWHSDNst87nSbq4xQzVr0Hj
p64HETmr3w6thy/myDDxVYNzoEALJGLEeQyMlZPnua6edEtkD/cfYrImthdKprUe
9HdB523zxNGnQIcAUH8XlcygtqLmJeUrrTJPKWDcnz9VQQ6NGfeFUm4YDXh1EM+m
AQvrgbs6Is8fzn5N5Nv4yolDJzLLYcDhPWTyu+7gFQE2D+WJa9Z/tpk/2KknHO/F
AOdd6KjO+XLk0n1ZQyt77jonzb+yOmd7FHc52+70NvAIYpJt9zkS2q+UvPhKJjej
F5cQCHCSQuEN6C9qsa+AXLXYIqcGTqBQyDLskASJa9OYgtv0DtT2w09V7QFvlx9D
MxJZbaXhwEYEjH9yu/JAouQZ5PEyZXZLfxLFgYETpfq5QUa0jENbcv0NU2Vk/EC4
LYCa3UEV/91yJh9hyP/0Kawx7M7xXUaaE7atg3jtwL/68pc1l3hgtsWZvRIlTpRa
tEDHctUtaRMHa5Tc4ZB27roqqgygL5m5FfpWYVPu5aPtSociG1XS+/QYEuvl8dXr
wYZfYyDbcddKQIXeaAx/kMGw6gqrtIPkKavafLF8PnIWs+y50WKo72eGX4MIm5HK
wn9TydswnDPF80cxVEF3DhyaqPLl5qm+kBgyWB2H3G6Z3Guzkc7i/NvGAAym/Bpb
vqx0mqZVgL8qICjnpVa/PaWj0QEbRUqxwnjlbXcmlOuLi0DFcJfyPtxSt18f/GBE
ydG89Sqwkqg7hYnK2mCKlnWr1Y8UHWX6wKMvxOccHpDFxfYUk3i5MxTR7fIKyGXS
56/Po8DPT0uhj4WUvSFCmILQB7B/HBIy11PMjoFJ0+d3EnV1VzN5QCx7ScfaKP3B
rhsMQ+INkHoTqhGxkx5YTtK26E5rYq5yd81ZA1baqPYSp1tU/BqzS3/8EUXEg2vw
gYmOei+EUwn6Y/ZkglpeTvsjhh5HTL98eKbJsPumjN+s7H+j3jNXoqkvuQjdE4Pk
hhuyYSh1yc5D7qM5QjbAI27W1eERHGfkpjTIG/1TL1h1pSJaxaxvLWdZ5XCZbZuQ
Qx7boUZBk7gGltjxvTDTxQVkwusK1tyS1Ha4QlTywHbdX3L8rOoZgeECeF4ed9lx
jb8T5vys5js4iFFiiLhzJc9rAvrtiZSE0xW8JnYNtlZ1pmli4xdUn5kGzG1ABPFp
ftgZ5wKzXgGgHqz1al9D5HAMHuWhEoCLxWW49N3IryAnoBNIGrdmas4SPT0xfDQt
xzC7GpT0KoXSq/8mTAEQL8pgO/4f0l1gsSklRkplFc44gZ3SS27KjcjMGGE1fHPC
jyoMhpkR9GrqRwkMf0xYVYCbVRCHLbzsFG5p/wMOmMD6cA3Y1Og2SIxmp3rOdItm
MnbxEA2eNHULeKupXVLTYsFWGGxoU6dRqCnOUkvC71zs2NnvlnYmGKl2yl29QJnz
ydLQW4ce0V8RBoYLsMy3w8GAkdnc/+SSKoVc6lrPM77YN0rq8angM6EMdNYoZLGi
ksE0huGk33R9Wx+KksKfG5p8dRozQr4EeUW6W4gxXKcgb/3Om9XGAEO90tf6QXeF
OhWJdG0REmj1zuzZuBApNkzKtSsur9YI06tYYap0lSbCx51x9LAdTYQPofhe33KS
9HN7UU6LBpNprPP0X6m9c+r98LjXcIWdKBkO7wzjDb7f/N+iQzriCFFy8EgmOXmg
HKr71V7JTs6ac4rJqxb23J21QZXzb9cA6yNFI6VuEnCCTJVcLs9ebnMEWOZHZIpL
MIOe5lY/dEKU3y1hg9qu+xktzRTIo+30UF1JsluSPxwUMjHZ3/YtphLaHB2KA3Xh
JnBzCqCaIED6gDkd9dS5IzyLg/WSzNOc4wbpQbq+LgE9YqgC69UfNLc/s1EvWWyT
H3k0AhRI+hCYa2Poj2sTdEbdw+WiGb04qD+t8UcJpFm+kkoywPf7y1vYB+Su7/1K
oK674zSp5qkr5UTHGVYM03lcBp/AChl2Hl7tFJVw7pQyMa76Qbjl2Q+pa9oDkvls
uX6HxJBdk1m1BNUC44YxJgTqOhMSnbs2I0k6lweyw8To740J99Dy0WqdXBEgTMix
FRUNrJVZp5fojkF5Oo6j5mUmrrVOWjwQ4jcbGRWfiBn2PNvu6Cs8AeKqnNY4Cgrm
DHW3TD9LiPb8E4QiUq0JwO1WOvDrzo2fZaiwgtpkQArkCSg27QtJg1lxYFQNa8zb
sCHmK/jZbsvE6dmZduNaoCxzJ5O1Kn0nDw4sk/vkRweWCnixorl1Wdt7Ob9usCmk
SMz2wPpyy1c06OOQbUDsWxkg7cT5Cwtj0er6t3e3oCmZBHiMm6Z6QNXJgOHOloca
LRAtlkdibI5A37PztSTGftH3OkjAnyh5huCTn5QfFHRGA4ZQWw3MDNQwBKBe32ES
CvpAR7s5r9V2KbGMdWXylZjCkHCuX2W1wRJJPf8m4e47ApsN8B4/Tg3eFbXSHejo
OGD6CZ11eXAfADWTx4FrsDQEo3rLnHM46JxhZt6R1x6wBdZ4cuCIjBSeFBVlhA/k
snaSXbHQrHoOAI6sOh3/8a3uscLd+lY01NBIxveDldLKN/u6PJjxYbxyRIqKEZgP
ADp6rbz6NnHzLOIIFQ7GLQVAd1j9wdwR41UkAVx59eETSpf8tOtYcZFAD7JAdKOJ
6yZj8eQwZEOaKr6imB2Fz7GSybFPFTp8Eb1JiF5Yu5sIO0vOHVrzcplGCg79mTth
rmpDlaT+dWS//z0pDf6ZdV6G7+du1Zc43j8W0qRNBhcYOr/WAJGJ7DGVNod1pIYi
rP9fd7lbCh4V2FZ9lHvg/eCoo76gvwp6sG0UMltJoAcTGN6QYgMYxk33OQNP4+Zm
W+XpUTrycIIqZYxinAsc5LsMfuVX9+VbZQdaoMWK4luiyGYdpw/vwr1zEt+h8sOB
BOcGIKu+XYgdeXc5U+Y+CWP5ostO9up2snyAhluxhgzNE0zIBuJH1/5BlBiQ4LFS
kEOwG/fgMOvFEbAhyDDS2dOzCw3EiP3YH5pnjRhx7QN0hocpv76485/8Av7lB7DC
5+DludbRA4/pgC/U+yw6CCoq5qxtrRmizQL79LWeSFg6tgBp1+fte+vrJa6d74Kp
7giKtmVB2GUooNs9wvXqUma3SZGPKZ2N2JFHjKxg5NgprQdO87RTwLdq71JQ6Few
UCuZ+dWOyp8tBllDsqugw8sxGoAqkdrdtrf7bdKmiSyxr+2GusafizcE22y2/9Hc
IKnu7qrR+/aXm3oTwcnws33kSYARccru8EnfSYL4kd+DEfTqqtpktW/Uin72rMhx
wvJxrcPzFZROnKXIvCR/UQtuQxMWapa8Mz3+HpxYUBdOPwZFG0WkdbVIRJ6bfMuV
4xdalJySi1Cvc0BfzK4niPSKsmZ7jAQigqP+2SNskVfaDdBczAjO7FbKUO6FjQ4q
m71YF2GfgQKkvkB9xuT80AVqFeXZtTs/QM7Dj8MEQVVASzKODegnpj/kU5rLImIa
isXyLHxArmWIR0gU6JxMLH30yxM78Uk/gsjEXyywp1CAS1227k6Ibc+YGPWdB/li
ps7ct1XStS+TIhk0h5bW/PJWtQcV6LLIea+taF8Do4b1hwa+6ep502afjUgGuYWU
gua/cyOgcZg0qd5PnFuEiYBijb+sVMW2SdV1/hka/FI+PXmnoZuSPUiTaj2ZS67x
hH/HyrAgsJDf/0/hTHK6eDd5cOgst9ycaI5NlhXNdD+gH5jomZKeKgV0dsWQeKoZ
N3dKjfzSuHWG2z0XpH/hb7cdYFqBhiWmObIC9sMcF2nURiRjNCernnxGoifr6H4M
leyZQ1jXK7Vv/MbV3jz+zNXCl79IawjNsufG2s8oZ0yYJhnlYoKJnvK3S39HUDBh
5EyTPRP4L+oh6UMmjhYI5pZd8iYopnpbB8iHKX8X+o7OwUSzjc7SRCJOz/VOvhal
4mJ/QNJOwz5fWqJ2HaVwD5KkmW08eM1OBgCXOmKXn0uWcJpyV9X5gqlHZ3ZXQX+z
a4DsmthqSEWic2Q3k9KiRMzQOUylCBNXbGycbMdra08F8zFhS9OjnQZL6xVh1D1m
jN7YtApqGr79U59KtibkQeVu7tTt4Eze6/nww6ZSw3XpQtoM5tHWkFmbgjdBDZnQ
Fp0nWpA9gE1Kv/RMnDNrepEqX7OK1+JbdLip5/AOL4sfn74s+m9+JbrnZ14iWgDj
+bguL9L67YlgCAs2l2ngWQ5ZYUHcxEYUU97V8rLYGEB41upyPWY+1ymy4mf8Jv3W
geexEAEZ/2FO1uHEZRKNk1Mxr9pRMn6ETohS/DUZWaXVd0VKRFUW0B0qmsyJSJ54
Za5BAXhzrxd9oZC8wPcdfSm2dBiLlzq7bSMmGugpppOmNuMkx6Sexlve75OWFJH3
FP05kvK6v48CmkHbjWc2Ds1ueos0gF+mgK7VH2StEXCq2hxmZIcAq9pPRMM1EXaG
hjaxVszAu/VPeTegtfHQgpIKP8Lqz20V/lOfN6GdUPYDM7+WORHFPznj2q0bgzMI
yA+CPLUgPx9G3QSeGoJvwCOrgGO34EqpKJflxumvHavKLPI3QY6Dq/Ixjj50jQVC
6OxMn3gzJYb3uKQ3SBNuFwDA2Mo8ri7n+5Au6pvR0I2dBE7PK2clPfX/IFzvgmLI
eZauztKxy5wfilCA2OnYJJUYusB9rZyGXYz7mTQtEy2jRjC6XbR4zBPxFylRcVg8
z7dxFHzGn5DJTzG1zR/FDY5SHxnFGSMxSupTmSNMHs3z18AabiqraQstxwg609+J
DvJZ4idhklFJlVP+6cgXtvzUzjHMxO2y9A3ORT0LQPpWHtc0W6CZmT4JW4xxPVPN
ONMLMUi589rd0XeOqPECrHrsZKChi9DrRermZcximumuylCInpxH+0XwrBfN5lJg
iOhYA1I9jxNECt6aX2fp3awH2zRUmbFJEpIGJZIg951T1kqq6yKFsw5fdrdMfLxC
0rWbZHAqHtBCfO1//H8k21WdfKzZAjwJMWtYP3Txz6iAeOshzQACzynh9Yybo43b
mSag+ATqspE/M025RV4cGcZLc31IRGVNyIghFzayEiZVj4//bnedpJlE9CIgsJtt
jgYCNnPL9ApX8yVqwv86XeT1AkZUn2trqqsNtgD8aYeh8BxwmeQ1ajU23xy8wYbP
cEQDZImUEzUTlhrx6nOGPHLX+/UjNlKHlq5tspmD+MPKxO/0tkGTSEqElQsLfc8Y
5vSNQnO+qmaBPQKTXExwO7scowk/MKzuKnjYwUKUqiWFNIViN+DcydWcG9EeN8v6
bBXvdCHNP5+prjjqy9hUQ/in3IKIh9zr2pLZ61xNcFuWgAylGfprS32DchaEX4NW
mHhT5gkV2leUOdKrFKajVhYfxB5ghLMk76Yx0AfWEaXwT47CSJAx4d68L5K611Ku
vTV7gMJQiRflNuKXjPSlTbf05HrfvgDPXFdYxdhwAThdgjixgvSopQ8b4Ljrdamp
xpYStb1JWVaE/EAautzteVHJeRiaRVmKraVak8054bxcSY2Up685KTrBV0IV+Wfl
/NfNLvgEqlZYoHXe+zG0T6I6q4pK4z+x8Uk4U0NKGwply7WjAlEJBYDgM+eB1Vjs
K9h9dJ31vmVMjYJQWBD5l6J6F/KpcHcRT/HN10WxnozVmLPN3Ea49niyicK/k3og
lIYiXK/EJjO/lwtXY3EQOilet571fwnyW2LAHnAcNLceLbFQoyoN5THotOSvyUqU
Nb1tGFNgTh2//e/BiD2QnMYldaoIarXqcZTUelYr3p1baqqwlY8xPB41pxVFlsv1
JIrl3Fbj/oI1Btcmga1aePzLW0i2gHHADqj21okjB0YL0zPn66sU0ZWzELuZvVND
WvkvM6G5Z137uJOn57+5Gn7787Y77ctHuzxLBgqSRqY69VCalOQGRd/nnhqqwcyD
YA/8anzfmSG81HCyUGJmJ2fsxIxTKu9DzgcAHi9WCTCvia4O9gcPOBaAyk5NGLsY
b8RzcmogObEZ4pAK9jSDozRfXtKMGEI+HXj3ReO60Sx/w/T/6Ieb1FU6ieHfNNaQ
Tk27yz3A5wiRz70xFok8Tj8q9NV7nGywoCW4aNJMnOe9n4Xq0G0tFr+7/J6vRb6u
KpdGVqny2a0FSlYaX3QQ3tOzOGv8GNEixcFPJLEe+KMyZh9SVOvN/yA6GNIrGxFF
Bi4uIUj0JrpWPDva0HElyJuTaHkBNP5N1A2TFZY5Zu/6jnGAIRxDbTCpqQe1AR6q
mu2gO/blMK8Sa3m4pi5Ts077jbENDZd0Y0gJeQcriItnjgLx7GR5/n3PKLCtrMfz
CoV2iDXUA9QSMVjpwKcFl2NmaH1Z5QIxGI/VqQSjHqAgrJz0mFbOlU3BE+5ZtF7v
b9OEcF2tDM0ZvS26aA9rwnoTx8xPonRRmGKUv52pQ8SMlZ0hEmq3QlKaT3NQQTPD
htwqoM4hOy42YZ5b12eTgjEWWQUOE02b7sLTn4EmmvjgOG1HPNTb1Lw36VSItLqI
kyXNlRBsenqtkpcV8PLfQ05EAi2O3VtOlNMT8STJo+82HYUg41Zq2Y6oVeg/Zwjb
Y1L7WzInJQiWIiw7u7YXCpBrLG0UaMoJHAUqvCNSlwcFcqAjyU9noYNaAmjQOUV2
Us9dBZQ2nOuFqf6dg3HSPcYdAKBMGLADHruqONmGOkQbXUnk/NlJoWeZK+svVJL7
DiO6sYsY+god1OboRgbQoNtrGaxEeJPYTlfL1m5kujObXE3F6SaT9+RjooaoZIrU
/Hwp2o0I20IfMib7bd8WPGYfODK3Bl/djiOE09VCYVZoQPFurkDiraHfEovNb3Yo
C947OnPlk4lrt+AfCXIRDkBPCE+t6uXHcAIttk6sXgE6IGAk8gPBxQ27WWY4GIem
agg+AHS0y8wFRBC1T9+XLhn8o2iYm88AgQ+PIx2oxsWBGPKKhJh3Tr9h9sa216ey
X4GcFsjynL30kolfPhJzDuswWc5U2rZU7LwnBP6WTuzlBJwLcOiuKsHMVhwsqiPD
XvOUzkCq8ulquW0KwiE2RLtAi2DjOtefYElJe9u/hm1zDulvVvz6ZwLucktdlO4m
BdkaDlvlbTu4xqHbgnTJLeCPEZCfie755Mm+wr/1uMspaQcJKBjZ1lZVpd0moNkg
jBqvMA450K/A2NKGPcaroRErqEKf7ZiLNQeE9FzzgyCzGY8AJ77NMSg5zbmMDDXS
XvwHd8mMLQ8jszNBVr8l7eo7FMn72QJ1T1kmCSDEfL+dH+X1lW/4nM2oKziQcqGs
XwNldSvUiraiUsZQFhD0mnGHS8CjrxRG38HU7ZsyISP2rFd62qraJNSKSFGYuT7y
ruC5fkzm2+AZYwHxvHD2wBTcao9NmCmy5EctyzHdk3/SLxCKE/CNNy+nZdWvYd10
irzFcf6OeO8hsnkgvPqAWl1VR2xoVYepUBiWHd2C81ZrfHEGV2BeJnFrFTDjpkcW
6euBYrP3fJ3uAq9XKtm2YdyLyPOfjfI07C33fLrsf4WKAeWWvG3ioRXg0TBeToQu
f9F7+RzNGT0fzLnurABb5URGI2pYhkFTFa5ukH+dVRIAvVqYbWo8J3vB2s7crIz9
0W7F18JlpTOPMuAHURL7bBuuYV1sC0BuIG/8pzFd4qTjj9HWLk8OKnfQ2HGsw5ka
0A0lb0veNgFKYPPTVkKSXBn4v7EiOMbkEKxkrxFvdktaITgCEzwq5CT4pEA29g/w
qFxcc4RSMVdCxyY+2IL5Y5n+g8+ovKHD5JRjDxapY/azaEVjq6IQwxwdZlcmPN5B
iI46MlgEsvV+T2L7MCNAmgqMgkvSO9a6m3EZxGL/ZlYKiCopI8GIgHyJAcDzt3PY
MsEq1GmnImiDJVn3GOhjB89A4DJHwQ9Wqw5B+brBCJP4jp7d/2JbO/QPX95Tvg2t
PMxIPUYmjYZDGwydoQTz7cw7dQBwWLJ9VKStSb1JYID4yl/fs+VaGF+3SZRKm2Xv
OheCcuzWGtFdgtkI4T3ZK5hGsEkOkFpTKS6tz8bzbxjWNtquY2sHt5SdBv/Mp/48
/lllRSV3Z8VXzkBfQEHgIhhpIblOoxFUFMSmt3QOz/L4ZfiqIctfTrx3Ya+BWYqJ
dLpqfXXRA25i1uZPjU79TSxwRtKCIQOhVIcXOU5znjMsAAGrlrzvcgjJtopeEtVz
Xw1SYbcMvngQF1g6/W9F7PVweQRNuwV0nkdDNSJRJLkj1y7NF/R6gmuaha5Of5Ba
YngWGqbg4DSJvi985P043ZZp5DDtxFULL0+MRW4yKiA8h5XWWmEbIi4D53i1Yr2A
EAfuMsVaeYxIplt9IZpYhmB7qGPQm5Q714Wp8eNBSp/BNliW1eDuknH5zLElNe0a
wvTrbDx10Kn/ztYhojubkijyeu2iqzFKHsFe5iN27QPzlwnwUEda03ATRRds+PBP
wa1V/SrcKPloWvTO9EXD/yujIkSkrAKbpf+s1KQXs9CTUpVsphj6FUa1156T8tir
667Vazk7Vwx2BEuPEM3WfShTjM3Lcmmg1HsUVbqsPCBd1lHYzu85rNJ1wj2yuM6o
kIIaptBsNOvxsLuSc+Jxw7KuBsI3WCLO96IrDw3T5bwOVqu1AN98E8foncHMSrAP
nJo4P8zmaEMPgkme6ZynCzhOLgglYwnWuVRjUMxiPDn3G2N2hBfMGJWcujCPl35q
IoBJ6hHA3+UBFP5kIMYIewbHxWoDgTL/xA4L/wUx2Norle4QiKmcW40i6mOFYfZN
7jPvHgBQUncWDjtUaA9dJd2S12BFZsXTFifdATUer4oHAKroSWyWFOM7udMUlBhj
4ylO2+xhnA8rA4v3JwSdVQ+CADwTqkerBVomuzsDRIAW7GGJdAulPGLfo2YhCsdI
o//Q0FuriSpWYqBFgq/n+1X8pmrDrBsSizafJpPw2mxvb0nrNq68jUjHJOpAJQ3l
SqxE/wuyHid2IjxlvcoOry3cLjsLyeABOnAqh/a45gpv5qpkDVR8ptIWcidkhkJm
ysq0X4zfaRK96F1VjsTGaDgGjnbVokPsIY0UIxsNeQ4SjBxHCTJpECU+zuZ75bfx
Ciek3ZtC08S6TMhCVSOrY+RDDUln9bMRcUD2zhrv0VvF0V+nQfMrtquUt5FCAL5Q
DtAIUg1t+Uo/BB3yuqHQoJhPbRqMPDGuosNhiWQHIT2uyrLTWwlqxukJ8t+tlpLa
gicaQxV5q0nPNUqhvf3P6TGck6mYGovq4tws/TiKwJTg3RPeTJHS1Qa6tLx61E8b
sQB0DVQDfREKgAiQorJxukvyP+s4d2eSKEDnsikNayoCAZDvBQstyJ/7QmMSx9OL
sVDR47MEBl9PgYz88b1AD/e8ij1mqTUScvbJrPkeMlbqFzpfHv4VFAeJV2uoPm3r
2WlPo7nAX3u4ZFW4Ia6/cwHtp2mPVgMqDxEgTpUo3BFmcc6Kf8x4SfXObeepPGP4
OVYM2+dF174assXOIdUudm8VZQ32J7GvMC5fV72vHPlDfNbywqZOn9jHjbZXX+f/
Iisf5jTAlw67AhtvmWPnL4EX8rX0asdjaF/FlI73p8aNyc9yqEugACidLbqy4+2l
+61B/zowQEWKYt/NA+Bnb7OEVyaTNRcZQfGwOxgWhMnQoRM3zdGeMs2PzlJdZyxV
zHx7S5nA05HsZhVkzCQ5JLPBFoo7y0tyBs+rYzqEmzyz0Wo/P0RtRHTlg64e0C/0
MYk1Llm2LE6M+8QQY/w4Yz3FMz9uQZ1z2SYLMx50GJRlnIQ2HSITg3XlC9S4M7V6
wKStYXHZhN6e5op8uK8L5FUAC0N9hmc/mSzhfmaNg/Hah141YNpbgi/3X6j3CeuN
JJngnfo1+H+DWOWmEVQf/IlbiSU/XB4mUc38btUvpergv1oAZ/6r2wO8FNJje7xq
bR95GWP7tTaP8zZ7x+bHun8DIQJYnVQODk89ssifJUpMBV3aNIj92VgAtveoB3Ab
zOB+Cd/bIUIKigsI5t/bWtoYKWG1dE81F2m4yRP60I3KknKUeN2wCwf/v6K3JDub
/JtkHg0g75cluU1dDOLyc2Z7ws2cZo1vo4go93rHlcGHBkRlcvwcxiDJ01eZwNFU
Nh5/P3w1EhNeJX5i3cs4J8HAH0xPhu+ON23xb5SDM+NarUwc1bOhA1id7NXZLovn
66R52fcp+FZFf9GvEGqfdRmLbGR2r1PTMnlQzRSCcZQEZhGBEs+VSOCXsyi4zpkB
Q01pRc2oANZlgBLzQeEQZa3Hb0Z8DynCHvn7ogbHrnxnxz36GnreTllfj/kwZEhU
EDJZDnO8oy4O7cYgKRuyuOtfXr+U4cbJ0acWTX2BVOow5U1bkbuu5TViXtdT7wVe
DfbD5uL7yROXGWL54Y/ZQghAX+OfJFdiNsnXZyYPc7xg3d437sVvK4AAJYD3nVDy
bU60zbcm4/wEC1q8EHsUbipArw+oc2wHnsiwpC/nBEUoH2RZrKVtUq+jHBJ6+CC9
p4Afua42q8+apc4KpwNfB9UhBIBwN0aZgQees90p51hRdgnH/Y0g7Wq7PErH0g6Z
rpp/Mlh3UkNIK7AetmRGE7DGdqK61ij+z7j5tuYjkVBBrGtA7CW8hxAhn1AhXeKw
GVw+24ngUphppK675zhRJz+aE9dR0zvP7BdjH0ngSSXyLViZRN/3nGv1TckTIItX
DswTEeFCWapDPGMdpipxyKK5VEgiYuhNt6KV9MqfYmuRfXldpS8ydY/h+1cKF9oy
N60P3iPcdNMshcHuIelEMLC3N+78YRqvIDtUXDQja+bIikhTumMbIt51Yjk+E0md
2Q10iUWWdH0/4en9U8J7hG2CzFBSEzrWiuaPuUyejQ/qlJKtL8J8ytMxJwPwlgtZ
lHhh4ct310VVar0ceiuuhScbkIavRKEplMMrNeL6Bc0v1TrI1pf6RvT7BvHxl2bX
FlpKVKDiEtwPbrFjQTt/mxrFZf7a8NTE2gr/wMLf2HwdB2m2N6dYDj1AhgPPANwg
jomiHGVXXUwSkjgEbaAgUQsaFmMXpn3UOXJh2pe5TcXhwNjxGlQYVSL6Xxi9obCY
J7En4yb+kZU5k9Iee/D9HRUAuJpY6c8xubS+5A7MwKh9T1de01exYPnX0dSmjaD1
haNtODIS+r7NP1YuLp+LPMNPFq/InNWK4GUi47bM2Hw9rSIOAMynoz1nuLYbIvQR
+mj9wUz3q72eMp7YyQzpj/KQ/94LS8bt9WnIZqjiAoHCQVYAl+NH0uks37yrFAyQ
OkGpJpmUxXarjjKxzDf70MG2tD2dA6JU251cPkHa784Ltlw6cXe8E1XCsEi82z0S
P9czmL1OJ4tQlxNEgEpMsmAKfN1PUmuOcWI0yzR2fVxXPeto4dMZ2vp3YmtSOiXq
PBRnKtUdzibGJuKM4CIZUJwkVeCmgWXNauZ7Vc61fRWPodCBf4DYUuHY+HHAxC4H
i2ofstDx62IYThE3fOl0kPyqGhySuoBz2n8QVkFW4VhOf854t6MQ5mZmd499sPpk
Ge6ehmUn8UEkARUmzOsG4vxFGRP+pNq0pibH+MP2b7wfnAOxjOr+taiKPB58UmhR
VU8A4f30eKWS9IyP5bFA37HKNBkLj4YkSD3NQABGXTMpclzr6YMvBwD4PZVzGuKb
N3wP9QCm01MufDiMX3LuwU0JXwcL3/3whM8H8LeeLd/0ZEtlp7WIxmcU68tx+fAq
K8JWlKDnR1T7ZuBV974DeJo8hyKKnoRE5Nc9OeTiz97DqQ45RVT+LwbIvv/FJ/qp
5HRJ0dvCghs8sjHouFerih/WnAUuvkIJn3K/4CxgXOXrWbqLjE9r0xo4LG0csd4u
Nctj5zWFi1P11aFvsRhnHKT5JnIgNyb1VdsZoVhnhHiHwzkyJMQD3W7HE12VFkCS
rCUMPESK8vVMA04NjOnkpw+Ke9qPIuT+1kN3sjEKu0YosDzRxjwWgQrNg7rkdDgn
Wkfbm1xrqeRUzVnNoWTgoUnqrF4sUeVRYTDEOxPzc07og49be9D2i/uEh8vtih/m
F8JhPdH5+j61BEeoHIBzDFUkiQs7kZrj9A9aiT9uwYvlwZPvD4bGsT+1AHm63o0w
yVtvLNap+MWRlH4wHN+LmjO9d0ATky2+lCQu/mPE29VaC2If2Gd6zjur1E7H8KUJ
NZm454dtOTxMuzvPEME7JSdMWhiSgJQ2rsVDqcb8MPFygvzM8+hbCAJm7p+3HQB1
vDMFBi4ghxkiratCE6YgmRI6zXRQPTqteP0P+7NvaPE6ocfxCciLzpSYoOd9FIkM
Os/E3IlU1rDwokv0xRxkzarh/NasN7scYfZf9BbBBHqJZ4fkAeMugDhzc29aqN8n
Wf84YRNudfRyuRE7C1aQR4esS1RsznmK5izBgrzRr/ycph6t7hTbHroGk7JcELn8
MlC4J6q6iVeNmROcPC7fqbzDkUafNWSRZJUKZ2QNs8YCExTiTkinlCwnrJddIipL
MFdpfB8qyINwffVxp4ww2tNGMHa19vTsFLKC1FHAIV/JD+03qtLRTCg9EePZmBuD
RM4fTRgh+qrWG7+7cm4J2CiiTYJcttPv0/uYbE3xcdsUi8LsU8d97JoqZoGdLQit
fegPu9dZOClA+vlTieGV/EBybH5FuqAb/1r5Xo7QH4vhpr1ySHOhFCxFJYN7dSUh
wpb4nzo2PHh+E5+zxME3w7vCLv4EqwIX2pbgQP5N2T+PAZXMYJ+DFEb/QFyku/sf
yFjioG75CxQyHyQjLMmc8vV5iV9x7GkIz9dAJ+Q7Dn4ePgHgGPDNLGsWdZTlyyCa
4Pwv4g8b6qro1krUlfCr9INv+fkVqRVnm8U+UJ3EkQj7Qw9Xy/uCHzD7XqxgiBPO
+bSh8z5jGSdGrQ6iZbv28bHg+2Pup3uJGd9G00F9IPskOPQ+pLW3ZbSGX4kM2pub
r576bXjkaTaDqq+a+0GLEyBsUVou5ADH8L222Jf4h22GdhVYUgETMc2+zMkEEF4d
EpXTnInCVvJpKLW0wrDXByElRcii8R/eVQ45+2nMym2tte57EDqAMmXF+4g/tvgB
K3tJ3Vo/u4rfYKp/s6EHg4nOJvEJFVqe+EYztZZfcFjWd+PAj57it7w2YdQdaj83
3CR/dK4tCrPdqoevUydrdhXExsjDVzneLEc8IDXiFQoX3mX+QFmX1FgIdErtHprH
rfbGLNTQZ4bZ4jCKIjXdxogL7iIgm7bBjq+RX5A5IOqOKoA7eWWf1gF6tS3kwsDJ
V9+f+GAd5PtgEbZpUw6LVmAvHEQnjyhZQSP7BkBmtsOMnXavdFtcsZxx/s9l5RJP
0T6vVYIkhShVJzoqVXCakEEt+Fe4gRbwj7IL1bNj4NUAnuTmh4jtvrnjcInNhY5w
elvI+P7Fpdc30yPG0lWVYeB+7rmLi0MXlV6VpXDPtKFDPSbuVrrcNvwkbLQeTmMJ
GvjCEKv+JW3yy0qIXILGRw/qrA8kIa/+1cE/BaNzroxNxmSINMJaCW3fXgIsJJsH
vM0dcAeuXKbdVYdxwcWhJ4wZ4pfnYBGsgBnrYUyVMDpqrXUuJEQXHhhc8XU5MMjN
3jf4oKZjrKKzULUnXn70mMGqRcPqfgqvVglCt0hIQWt7sw/mf4qbXrpLogaMeAK4
Wxcg7a0RMqoPENzXexc5WvZRw9bY/y2E7BtmdXdznQH/iSoP0CXGHwiKGj5pA3HQ
8FSkcyyjFBrcm6yBIbgf44I9DSD1BKCN7UhhXP2Ml5CGDoOzm/KR5cKafVYj6Oe+
0DcLouhIBEgfczJB46b8Lc81gSZqD1+9BNyhzaZVwtZuAHMfmT/0y0X49VSy26PI
//pragma protect end_data_block
//pragma protect digest_block
yHWvlb/wS1VkGkPXRXFBErSdQ3Y=
//pragma protect end_digest_block
//pragma protect end_protected
